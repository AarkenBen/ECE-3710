XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5�o�%�g�-û����tz���?�.�\��G@].Mg�'����"m8Pc��5��9~>�*f�7�����ј6���xYl����Ec�,év���R�"���<X�'Na*�l���g1&B0VFݍK0����a�Y�3?kSMS�$2�����L<򵭼�5��J��I��Ӧ�:�#����%�*-U�ڻ�]��FTV��ش�Y��c]�٦ϴ���S4QV�=^4����
)�/�����/�Q��z{Q� ѷ�z���� N�/M[����o�ʉ�v}r��'��ve�υ��y�{��Sa_���tI�I_w��%U�O��<���a���}����R]&�F���"���|�y�S|�H���n� �e�,��]֫�Qa�2��Ep��O�p,�]˾_�R�	�t>I:���9�X�<8>��kb�-�������R��-��CGMp
ԢWaM�uS���l��J���v�~��n^Of$���15?ࢻj- |�}c�6����"�W[ډi�k*���c�R�՞pCg2�x���kG'�� H>7m�S�P�:w�
p�i�	|8D�:����X[씪E,1sOWt�ͣްmA��^�����{�x��W�)[|�w�)#6�cu��bQ~�e�Ȥjn�u	�'�3�GN���du1�2�.t���֯��w]#�p�q��a�� ���^K��B�	[qm�6) �m�a<9��9��gP�`��;k��t7�����OJT*�դr�XlxVHYEB    fa00    1790p�MЗ��)Z���ѥ���֢}�:��e���Q\#�e,����?҄�݄�bQڮgQ%�R�U*�ܩ���ůh�6��W�
�^]��Oi��+�6���g�����F ��y6�Z��L�F��}]q���K���hp�o��hf5�b�U�9�㐉��^�U~~�l�%�{T�R�s(�V������v4���a�g����+�Ө���� 0ЈT~{H	���!-η�}Am饴f+w�HAkoo0J�� /�G��0���xvN�`9�z�S|�R���(˓��vN��Ts� G��Ld$GŽ��p»�h��I�f�2ӗZ2�3��4P��\��=r̹�A�1WI�a?��C�m2�E�r��;=ܐ�F�M�U^�B�!���f2�uSO� �]�,���%�w4�w
��E<�������AV��51Q�X����53"Z���wۚS'w~���7$��.���@����OI:^�����"ǰ�O�<G���}},g��:�`��5����������E�_I{��vW'ō�\���-T�C`�"R�ڹ��c��v��sE�b�!AZM�d�%|�ϓ�8ɧR��Yn�C�
����Z�~'rꋧ-���$�y��>E=z�|'�11�>а5�0�}�������<af�/��2���Wק�g��GB5��s��T�qS�c
�|���Ԃ#;ZO�7��-r�j���m%P��p��j�M�����Ix�!�T5@���U���#Q��3�KL�ϱk�Q5�O��b��8��/�IzY���p#,���
�6�Y�Ve���L�R��g独e�������1EV�3�L�v ����C�Nw����s����?�Vd8�BI���mb�˯��v!����_4�
�;X��Y�ft���c��
��gD�Bf�[�Sˋ��f���)"N��>7v�!v��S�����Vso!"��.h4�u���$��e�	o�콎F)�>�+�MFM>d3د�����J��V:���R75y�0��)����Ue��y��8��^������|�j�`��ϛ���w�Cz$o��S�F� ��,z;�������N�U:�.�&G���
��s�Z���W�����"��v�FX�~Z��omx��������h�;��0Ef�չ���*oXAD�t���BU�_9��h��o��	�������D
U�����~u�0�����٤G0s���Ưz2}���&����/����[L-��@��� T�b�Y7����._pJ������Lܫn�.pu��d���˪-myYr�ӽ��_���x�O�㸉�%Ԃ�����x;��MF�����_��W�{�t�<��
�����֨�@�m��,B��R�2c�Ш��3���7�peeG����療����]��,TuB���f�k�,��!D��1GI^m����YW�3�$%
	U�U� 0��o�l�Y4�|�K��%T��5��[+�lQ��I��L�0鵤����'n�)��	/�?����+�F)D��f-�n��2�+i] ���&N`{��q8��2U����S�6����#eӷf�Q4����Z
�!�:��3diG�!r�՞�S������2_Z��A+i�,�R8��$g�����p�ݒ���:�i�KN�l�����55�8g�M��}���'T�E ���}e�ޙ#<�E ��d�^�Z��y�wBg�j�����\��z��x�
Wm�O\vU�?ܴb�������~�Ie0�aq��&��9�9���PB	�������lx(p��f�R��s�d��0�] �K�.��e�f���!y��,���I��a�bwѥ��m�%P/��R�d���R����!g��G1���.e�($�p�L�m����'��*�{�r�i���_���.���qp��Wn=l��l�dSd\�f�t�{�}�T� g+��RW��:��:�KF�J�9�):jݓ����پy�BU��4�J����gR4��	�-*��NN�Ŀcs>�*��9�g�h
��C9;�g2�T����k��O�e0���(��g�0'�*��	��%�}6v �#�ZpJ@�o/��a��yY��@�dd1Uf�Ϧ��� ��R���Ļ<�A�`��QTn�h�)�:) ��m3�������5����z��)��.��Zk�Uд�Ut��Å|��l\��g�Ҕ�ʳ�R� �@jV���}e�(�1d��ܯ�z�,~{ǥt����M@�_Jn+�P��<���pGS����I�z�[���dܒ��|G��}�}��'K2.T-w$����!�NC���F�0c{��m������]%�J�Ĺg�aw�Q�SB��8���@p��&jV�T�dOPXV�Q.�{
'���n��2�/kh�������|����Y,	��C(�i����:&W}�[��f/���m6X�ƙ1�h'�{15��	�Ј��_B�]�-Q�,��3��D���/�F�0� ��;�F������)n�����H�2!s���9�r"�_yD��y1/H�Z�7�snyk���ӵW�Y��'�q�_����"�|	�#QJ��q0Ɓ�A���p�q}���,h�T�՗���a�2!�q��Ka�OóJIsV�V���@�_�L3Sk ��x��tIT�uN��Xl���f~��H�a�Q�EvQ4��+͝,Ph*�a����� ���lFLgW��
\4�Sp�l;�#��A���UN�XW؊e��@�8��Ի������g�I������@:;w=?�G_�<{�����NkT�\Kג�������i�,�D9. jW��|����b��#���,�hϦ�m�xA����e�ιw��Äm��Zu�������f�|�(�щ����2�Ls%��S�q��f�~eW��4}ݝ���)4�|(��sf�����9�y�x[�$�/�+������:x�WK��:��.��t��m�`i@!�K�lyӴ�����$V�b|Ot{-���B��!�e"��j����'Lm�0V(Wy��h�['�/`{�NGo6I��ݘan5c��EdC���Smm��'m�Pjɪo����h�X�ߪ1`�<�������� �*ڝ)�!F[u+<�')��_��uK[]F�sB孼�"12L/Q�}&@Fv�"aS�$Ś@����8n�%z�܏�5���,^��k��wz�/d<�hcar<`��g@����,�a�6ǘ���<�׶�w`W��`^���w�@1����t.� d�����U���e+Xc!n["�|��G�����@�>�n���&dpK��p2K��������vAQ\@��=����k��D| OaxV���~fZ�P�)m��Y�y\y�	�Cޱ�p�jo�&� -Wxm��&���\|�C��kh�<��!<"W�
x<X��L0��#���{��]��۞w"MY�V�{
��<��'��5/�9�FQ��nO�δ�\�2W8�]�8c+y�9�4�8�+�]�w* Ǻ�U��1�e�{�|�3�m;Z)C���+�?�<���.��׳�$�R*��Q^�[�Ù�[��8i����]X�1'X*�m�5&�-Ƒ�/��+5�3�jn��ڦ�<�n��9M�ۑ9_d��N��!�d��W(q�~Vq�%���"��Jh�&�����*z���	Q��* Ě<��As""q�"�`��-��"Y�𢚴��LS���H�AU���L�ʨ��;K� ݜ�Z���L�ȉ�� �!���;�⅁�0k�f�'`���y�<,Mځ9fQ�p_⥋+�6�0bd2��&Y��E,I�m�u8��#�U�\K���"�Oz&U(��Jvk~���vƓ��<Ҽ�H����B�����/D*���]�Fk���ס��q��ן����U[����JD����QO��7M(M��	\��A[9$TF���x,�Q��
��
?鞽#��|�3�ܪ���IS7���j�敺��:�~���d������d���牰����Z��H���1�8�U����oW��L�<�ƥՂ��+"���{��0���!����&ġ��U�1�L������]/؍1V��ԥ�~�����៞gU%W�j�Z��*��	ex��ܑ�Xb 1�	#�����D/s �t�����d9�o��!.��"M�ʰ�D��V���M��*ی|0=bE࿑��	Y�ܳ�.ڝY<.�������e�)�%a���)��~�c��e�s�g&�)m����L6 ӡ�k9r���RW�l�Є�9��]��M�{�����`�f���dwR�:-�����o:E�۴k�@E!�����V���<��=r����%A���V��2�C��#1�^���d��`��\�G�#:Z��:��p+��S�b���H?�쵝~.��-��j�^��q)�R�dx��	�N�'?�3yš�
�n	q	�[�?�,�m����`:�ϋ� ��S�[d��g�ʤ�Yp�a�(9����.~~	�PEl�)i܍;���ׇ��9�<Q�D`v�wARǐ���)��{Bgq�A�, �V2�4 �[Y�.��sF���h^rB��#���>���9��Ԇ���a�]^b���d��@wdb;��Ɛ0KKu;����R1t�qX*z<�Ҋ��!y�����r��FةjN��k���\��P���}�P�g9t���Z��r�QXn`L2���ĥ��ɩ��܊�]�V�g�g����;�Pt ���~��Z��8$YV0� �!���6dW6�.���������L9e���[@}bga	Y9�f�� ky��ؕ�{e۾O�0�]�������z�?�~&����ڬ$p}���?�0��м-b�veX�K�����-�kN��s�]�7,`H�BI��	��I�X�s���snj�-����A���ʆ�ט��0f��3*����Ne��/�3u�%qVG���f����9"�M^6J�ݶ��Q5�?��	��B"�ж��\[	��ۺ� ۾
��h�3����}d�=�R�c"5B�)��%0y�u���o]E��M;B���f�װI�G����$���
�c߬�,y�y����B炼s���B�ǜ�>>��Lz�tO��U�hz�z[@��{�#��ώ]j��|,�8������z�m8mjECk�D��4\ZԞ#/���T�
5�0Vy�4<��>�Hy�h����Y�|���^��.f��Dk��� 0�T���E@x�V`Rzt�#bGq�$����������KNf��)���D`��v$�	�Q���v���B�&���8�J�> B<$�Z��:=��x��)��u��4��4��i�#cJ}Jހ�,[^F* � K��0�jE�9&�"�|J�c׸���
�J�F�A�žX��%�2d��0ʔ�����*r���A6�# @i{q��撑	��?��>����
.y땉��?��~�Ƹ(��<7�1 �_0�s���d�u��-5�v������=Q�K�Q5_�:��C��t�p�����x��B�Ɠ����yE��,�y���O���ן��j.�@+���0>��:�=��^ʓ��t A����.��O���!�Y��绠9��T*�%hP&y��/����#g��R6C��hw�:�������O/��QIr��n������i��C���W�.ȺV�Ւ�(���@�6�X,s�sD[˜��8�j����?��OQ�>=�����3���#�<�g�������S*���-��](\�E��h~b�t�ڿ�L�{J�J��M(����rc�e��ϋM�E`��o�U��i�zm��~�l>���;�aEIz��4?o��C��fh����=e�v
�G�e	o��f�?_V!#�15���k0�5�`oäAX��fS�#^�u��r��TfB0XlxVHYEB    fa00     5d0>�O�[�鱻�t	����5I��ō4VI9�_Y~�eҌ!-Z�8��oq��$�~��-����ŌRbu��%���M�uN��.��oYS&��6��P�e��Fz'o�� 6rtP1�Bͦ����ud )RL�9�L�����"��ε���~^uЋ#8�
K�1����
J��VB�c��a�L/�8������*=�y[!�ϳ�&��|�8��,sW��P2K"��~$��Zmóc��`�ՙ|�i�ׂ�{v�χۘ�t�	� ��RE?��1�6ԋ�n�d�ak��s��܆[��`V��S�Kr��O� ׼��/W#Ь�K�(�U2~S��*x�G�����S_:5m�v��t)bװ�m�Y��I}��3/�1� �j�L�]^��L�Dp��O���vs�`�̯?���(����Դ~�_�_��GL$�8v�GC��)������v[9�:�A~�[����]�ގ$B��(�Ɩ󾾎q$��
�@rj����:�E/D�	�؜h_�#��)�
=��zf��?�\����!��E��,Z�f��3{zb,>�5��8�ˬ"<!���9�t���Y;�`�͌��Eh QS"#)�Т�!�O�r��:���	���N5����iie��<�Ϋ�L[�e��f��(�`�Yp��/ؒkK<�N���ĝ���c�AbJ��US�J��9ΑR�/�Z���b�n]@�Y�D���+��;q߼�~�-�.4B̟����� 2���q��Ҿ`�?pm�N,�*6�<Օ�,��s���I͜ �G@��_�&�*T�6���70>Î��/����ϐD��S�qS�[~5_W]�~�xv_@�����d�v��/����F�T����x��bჱ
|S�I�)���^��F�Z�C��$^�1C�K/8���/�D��Nn�1�3�x�YSwR��))lO���Z&���7и՗Ј1,tǋ����6�e�,r�\��?}CY��Qr���glB�w$J�!6O�$�,�D���R(YƔ�F�����Y{4:8��`r��[n�3ZN#)�p'/�����x�7e�c���>�5���>/�������3�t�6s�$-i�J�O�k157$�o���]��lQ���y��CG@�t��WL��aaS�	V.����F��(�D��%TZ��ԔF���w�")B:�n�Sep>�̫��z��QQ@E�z�x��`mN9
����_OGࡓc�m�bҮx�mԓq���3G�������1Y-/�ψ��ҕ����/��K�m7-�tp���t}l���\� 0�.p� �}��4��*��p�*���tF�����{N��l�+��I#��!�[l�.�ȸZE�^p�+u_��+っL�"o%RI�V���جF�K��]^��Cu��h�#3 �ɑԁI��2�0�w���TKΰ��� >�'�d�6x7�!�|Mx�@����K'�XlxVHYEB    fa00     640���}�d͎��g~}��&�,{"*���N^��z[ʌ���/A�X�_H�%��j�B-'ln��7ҎU-s«��+��SKɣ<fQ�
d~�ā��a���䧣.L�[�!G��,�~d����V���^�@Q���@OϷ�P�u�����������q0��a^�V;�g�A]��i[o�L1�$�14a�4`��*���1��>��T��� >��ו���M�*��e�I ���Ds�e��ЇȪL�5q<�4t���SNy���q��-�M'�0Sk���O*��2�e�k<�!�jӸc�H��E$�u���!��_pr��]�����^�܂��gLk�٤��a<z�=7���3%K�]Q�゘Wa�Ճ��eN]]�w����vi^�+u�U�O-�2�Ʒe{����!��y������b�x�x!��E�4��	i4�~>�&R��g��Z��@w-
����sĦ��[ן� �W���+�s3&���������A�����b&�����ᮡ:E��V�:5�4�z�C4�h4Q�j��h�Ϗ��42����F6������@ݗ*�}��2�2��p
���F]�ܽ��1����lҾv��Ϧ?)����������3S	�4L����@����A�w�%�t��&�(#�K�j'��T�T�Klw�ɯ��B	"N��{���%}7��N���S6bbaZ��U��7Y[�/M�ʬ=K��B���Ѡ���q�H�/UO��b�z&{�_���*��;�.�\�Xo��F���-�g�WYxI�]x��[\�{��O�Tn���R���Sɸ�@�6(e�Xվ�9�d�Ϧ��W�Qb*v#�{Ѥ�u���PX2�emn	.�*犗�RxwK�+X��ld3\p�g�=w]_�*�h��}�@���ӌ(�]�C��<픡䦸O6/�.��[�Z_�` r�l=�y� {�ܻ���yKV����֧�5���Y�z�Zk7A8��yt�ϲZ&#�Kdmq�f��wȱ��6 \@���8���?�R���X�i9^��:Ę< z�-�D�r�hz~-�`�k�1L�S�41�*����*�_��w��GaQ�m�8��pZ�+k�:�$'6�>�ݤ��k��h]Vz>�6$�0����̪/ 2Ek�߇�	�r5�鯅�PΠ���@�m�L�%h�P�r���t!�YN��}������ȟ�Hf��k*��_���#7:���Ne���(�)���V�����i��"����ƜqW�ʈ��E�Lm'������#HofS��'�96�iIڔ���{4�{ f�7(	!*��,Ixf�tHM�z� �l���}���*�x��\p0)�5tI, �vw� 7���IZ���R$��m�������6�M�_�nA�b�lY�<��z�O`�c�x�P�����Ƌ=��
%��;��h��\72>�0Uh"��(	H�]��ލ֑�;���.�FR�6�7t4�񔨬X�p�$4ʣ��el0�8e���M�]�Y��#{"E�VW�ɟ1W��β�B���2Z�,�4r*`/�*# ���/F���GH�r[Z��o7�҃X�>u'�4���@�XlxVHYEB    fa00     5c0�
�w�U�7��TB�'��,8�����8O����Pn��opγ���n���C�h�����]�`6�OȮ;�*���껆���ܨ�)�9�X�6���%_���p��Yq���岓1�=O��o��˭��t��2Ǥ`�a�&{D-y�fg���z3F�DoSX�Z?bh�e�E4�i�p	�-�P]!�R8���/U!�/�!|r���Ž��W�W��V:@J�zJ����)7͗�ҕǍE{�d�\t;E����3(�jfW��������xL���~�so������5U3��[:�<��fvp�:�=j@�V�g�8�㽍/'P��BC-�����)��K"J)��b�x�e���c9p�[[��9P�<+��K�v=�Q����{Yx�'�ZQı��u派yfmd�_:��䚷����Zs�L0Z@&p<�`� ��ݲ<}�Ń���,^+zz�!O���(���@m��`��<y��C�����H�O3CXȹ]�$?�0M�<��ܲob�օ�ϛ��/Y ���ճ�\��k��I�l����k�hm�l��ܠ�a�˕H:��5��Y��C�#��_�&
�M��f�h<=V1"���x�B�B����QJ������꧜�T�7��I��t�c5{�W�gۑ��?o,3>�o��H�x��' 3h�����$�ތl�o��`ɋ3~�y�O.I8�:�u{�7�7��.�$wJ��}��;6�*���dA��0����FV�*[�~���7���cK�����H�C�VVj����^�#�7p 6@>�������ty���(��8'q���"�z3|
�u�����Fe}]��L	�3��8��u8	DЪ�j�1�8cF�e�D�� B�M��. � �Ֆ#�q���L4F�D�u�qw��Xv�~��B)RZ��T����j���IZ&-����.0b��ٻ�ğ�JM�I�Y�^����ޘ���$���8��T�q4�����Ņ��<�\�i�g���υ#��*�g�̴T+��y9M&y�uo�|���R+��z�@��T ]�p�a�5Qj��.V����*Лę�R{��':-}��� &ūOu���T�R� '67�f	����b�n��s��f�bş��?� ?� De��I-�."�C�^�>$��<�Gr�m��W߽W�9��W�I�oD��|]o<D֛����P/��ic��K�(:ʀX18�P�z���l �UI���+�_��7��_�h���D������dخ��'�襖���Z��c2�a��*�E��<��Fd�tf�ۄjp��Y��T��_��z���a+M���dIʰ�q�{��)��2��G����ܚ�+�*���|�{+C��7<���EGt�0�����˦�-Ý�d�ku��6��ɻx�J &�7�������m
����3���g�x'�f�w����/k ���,�j6�,XlxVHYEB    d347     a90�`z�pu��UI�O��4�xQ9k������Q#����3�7�*�"� ��6A���O/)1��j3�6:�ڍ�m�W�7�F=���s�����殒���\R�IqMH��B�0sz�A]S5�L��Yr҃��.W�������)�?)+����ɉ����M�0b��f	4�����<����R��@渻�f�T���]2*_�~	�� E�a$��e��=���#��b���{�;����ˮ�-Z��W��[]��!M�������Ք4�5ѳ�ȕE#���\ST���b1~P���`�NW�H�V�D�C>�J�دePJ$�T��p��uz���锁�1a�vKzT�������N��-���fٙ�K�� �>e��wf�$�G�g 6(�r\�Lйo�bm��R�;��˲�߬��0�}Q�X�0t�ء�`cwal�������,\s�t�#w/N5	s�nMxA�{P$�|쇟.T��Ăb�f9>}�e9Yx:] ��BI�'�!N�x�I3�=�r%x�Z�N*�������?�"^"�t%r����5J{yYg�3�p
�����n�0.i����7L�(���|�d�li|zAQ���-[�R���t!F4�,~�;.����l1�Y*C�YЍ������CC�U+���E�u�d�E[����ӡ��x��C�.�d�#��>;V�H
:�J�{��
���7{ep�g�Е����zs�������#�R�p��M���	*����%,�̸�4h:���+����	�yZ8�/A���@$�}���
r��ˀ</I�I4T�
��6����٤6-�o�ʹ�8�(�#\ى�I�nI5�?OS�&�#̞)�<B����!���n������"?��/uL4��^SC�۞z�Ì2���D��Xng�PG$]a�V2݇��5"oa'���(��:� ��:�?��ݙ��4����ͺ�N����W
f����Y�{���e��l~�H"\
3�JV/Nz��C.�5�ғCd���&m���`n!�]�B�_}D���^�uK����6���*�qe���!����g��@���U{�@��W������/�w�rE��S|�x �3����yJ�����D�~�D.�����Jm L�v��2Ϟ���/w�S�~���@!!��Ob���jhDܶ+�>@�x��*�L����є��&\�����\�L�nb��~�/|����{��"��eh���X�fm=t%� h�}^(�@=�YKA���%30���,e�\ܙ�k�����s�G�F衁�m����@��Z�Cb�s�b�]��hcH	�P�&	�|`��ܶ��=#7AC�f+--%�8��sm��q�wg��d�"Wj���a-�Z�H.h'��C�{�4�_��Zx�=�,j��b�˒�s���":�o�[�թVLY~��?�Rd���I|�M}u�li������sW�����[I�uk�d���!�)"w��NxN[���P\�b���B̈Z@�[Xpc����̅��<���|0�3� vo�`C�xb�6�m��PL4�g�Ԟ����U���v���>&�ұ�l�br�1��4�J�7K�WZ�ZZ���B6�D��(qP�hka���ߝ��w3q`�sƥ;�9�U��Gw&E�E���j+��|kle���لp�Ar!?*�F;&���/�[u�e����{m�M>���:�I-�g�PyQ�3���0��0��3_�geO�sB>R���H&��@#��1� 0��M#���{���p��O�y��/@@�t�`.���.���p�5?���f�i�E�E313W��$r0�2��my�P@?�H�F��xso�ij�u������ )��>��������1���QE"�3�А�qR��i����Ж R%գ|����%8�1/�Wv�Gr���kN�~�v�=��g�����o��)J���4U���wa6�PkR�< O�R��;u�|��Oq���'��f�3�d� Y�-;�R���o=k)�����,��I)�}�uVkL�3�J�K~2٧�p���eN>>	��=�F^�����,�YiG@-�:�Ռ���W�6[�vo�����9�yi��G
��,D��^$���c)V�zW�-�ߴSRN�-
�aH-�2�">����+��rdUξ�V��TaZ�+ .�ql��c��B��ޝL�{@t"����P�h���G��Nm�N��~�ӣ�}k~��1���J���`��Tj`�[)�eYL�:�Y^��� 'U��&��?y9)�fk��t���.�o���s���/i]
��րU��&�а`6fR��raf���$:]Nu��̆��T՚�,x_C�֎^׷]=�wZ�� �~��H5�)}�i�f�[��v���s�ȅ��S��� �VqT
�J�s��/�wH��L�uŅ9b�L��:�t�y--i�+9xdD�\�pwO�q�0X�m23�ԍ�Q[g�O�r��k��xG�O����p�����޺T�����/�C��d�J���P�4+|�x�^j��O���`�)�|��}�JY�X�e�Ҁ��P�2�T�-o��U�ly�귇���!��rFL�dh](f��U���cr6n���jW�A�� �U�L���ݓ�o7���*�)�����q8��