XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$	y���%V0s�ag9�.��q0���+��Q�a��״&�dޔ���A�氘�љ�"�t�i7��{}�3 �������Jx��������[��7�u��Kܑp,�S��&��-�g�o��ǰ�;+wgL�Q��!q�3F�Qt���}q�����"I8a�!�1rW~��7�&�^RF���lL��@b{�þ�B�����8��j=M��&�lk)P �P� ���5��nU�ůR�
mw-�#��&�R�]�6U,#��J� �j��S���袷� �˪�A������m
��GO���@���fi2x)��;Dm��j/ы����"�&�pA��Ж˸�I�EO��&�5�'S.ս���~�x� *U�g�����.*S�g�/��!u#�ו-���$C_A3jm��N�t�\M�bmS�I���4�����5�)��d��:ym��_̤"I��W�)U����I*RŹ��_��KNIp��M��铆�-}�&x�ťzt�N&�]nX��Ne�ARu��F�"3܃%S�@Ryۣm�W�6�7"uS(�/�s�� X���G;))H��ۋ"o��bμ������:�k��#̿3�T��8ز�4O���.��6_���V�-�iA�iۀٜ�h*G�������P9���"�i!��XSҧl:=��b��͇�B��S�Oz+��_��C�2,�m�%����j6N��bڻ�k�͕� �Vũ�Sx�����bUnI`x|���F�h���5X��XlxVHYEB    fa00    28c0YS̙6<�U�o��]�zڨ(}�����&	�ag�O�XGc��6A1N��������ί	)tqu�jy��>Upu�+_pR�$6���o$��b][�tIU�7�y��J�mƘ��O�:7juݯG��[�ʙD�����a�I`��}�� P��c�����r�/_�2m2|�	�H�٨~!���FJ#��*h?�J^�B��@�I|8��B�\>�/ �K��j��E~���"��iq
���=�N��rٌCB���
�= �G��?o2����#��m��Kl{����FC�_���nBٌ�ɘ�*�=�8�λ�(�C2�d� �A��;yjh��.r�����ڲ������ ����ƸE��i2�8����`?*e�ABb_�
� ��y�;��Ȏ�l��ZY .�:(Y��:Z8M��5Fl�U�z�F/�ǳwZꌥ=���c�/�^�#ɴ[�*� Z;�v!
Ga�mI���n�^p��oV��-{������5.4[ ��ڄBۭ������5� b3�8-ŋ4X���f�v���7h�ޛ�$��A�G5�f�u(��$�&5Ӟ���)������0�R�-���y6Gr���=�Dt"P�e\��� $�=a4��I��~�� ;^44�O�A��K���!7�W�$�|[�Q�/�J���;��%K[��pnO�� :����$��ۛt�b���<A.�<�wE����(
�!\�Zٖ�3|D���b郾�N��K�����F�qZ���m4��~�#R�/!�-���f��a��M^ɚ�h�_^qˢ�hFU!�@
��h�����)�Y%@?�(Jj�BXQ2�2�7}D��AƓ�Jj&����ش�v�+�:���7����[N���l��2�
�V�� w����42o!SW���*d��kOK�5�}���j��8տlf�Ϲ�p�k�:��Od��:{��Q?ZK��L��\q������� �-�$0kV�N;%V�*0|��4���u�_{�/{���̎���)���/6��qu`�
�Z���4�gKz	B�?1����{��(%J;~���>좸��W�孂{�h��x	��X� ��.d��/	����RT(��*������g��sQ��޽g�ˆ5�.}����\��GQ2��A��K��A�oz%�Je�'��:;�%-y/���1�n�=oG��ʀR��2�@��gA�Ǥ��!�A��aT�i�O(Q��+�GAx$�K�4e(�I�D�8R�+�h����kDK�������]��k�<`x�����^5JmWy�mS/��e�(���BkęE�&�*熲�& O����L9�����zQ���Q��(Nx�,�"�x/�H��֟:OL/�\�0tMj�왱M���U��n�x��쥥u�nR��)#'\�_�ך$.iz������p���Ċz6��G9n�}W�V�m�nBX���֙��a�?o�]��QM���	o��B ,�]�8�g�pJB&S�T���bD�D�zrN��┾5,[h��)���8��[ɏ��(�xӮ���!�H�o4Z)�����0c�n��T"�� �J˫-�BAJ+��=�
���]ް�-m���|cx?��UCptv�-~�?I{Ԇ�����myM�N�,]㤧�@D5O����>	0{wO0\M\�Nf��J��^l�b�3@_-8��'�a�+�T��Ԁ 1�]{s�b9M�yn�*�ȋUH�¹�,��Fޠ)�v�q&���$�������n�1�_���;(�\Ir�s��$zN�A�����	x���v�T�!���xN���u�Z�P�v^8"���<x�7�\��
���\"T�f� \�
1��T�4�J?O/��jL�)��ӊ��<E�Y&�Ms��U_���b��3�Ϛ �D�>h�+��(�L��J�` X2>@]%;q9����M1��,��(���.���������᫠�� ,���ֹ�$���6i�ϔ�p�Kϖ�Ȼ���N97�+J:�ȀP�?c&VaVm\Ċ�Wj� �ϻ�c��ݩ=*�,dV�bcM����_a�*ؗ��å�����),�;�OD�<%�V��*�����87j5^ �6����M-��y��/�0{��9�!Y��!�����Z�E(�݃{b�Ђ�~�BpJ�����'����L��c}�=�xaУ#���N����;���Wt�
�[3��c+56��	�%ni!�IWN��@gI-��H�e'B������(�Қ���l��l�B��^+��U#��5����K���<�0����,#.�Yhi�Yge�E!C�<��1���7�qV�w��GU���t5���������4"蓣��
7q�wu�� nd����s���d鞱�m�S�Vߘ
^�+ԇA��wB�N�eP�?�<8���p�����L�՛,K w[�х��DP� ���`=4w��v�j7ĕ�=8	�V.��-t~nv��FxC�тSm�#���2`�c���kA��ݧX�W�]X\KPH���Vk���{�֠����:����
#�C�t"�D�/�30�)5	X�r^��{f3kFSF�0��sG�Q�@�}��UA-����EN�\��D�C����z�Hp���������r���}9&C�(Y�칤�B�O}�!�<x����U�Պ'�E��.���_�n\�F���i���%_���S��Az�H��p�����ȯq��YUK��O�z��u��kR�_s}aT�NHⵊ��{����0#�6��w���lp����Q�l�~��^�!������&�	�s:���_�7�Oλ��b�V�]�1s�"R����C
A��Ѿ���㤞�
ݓJ�f;A�e-��x6ueృ�p�DW���9CK\ѥݭ���Du����}ڶ���PK���fV��l�~�+R��%.��k�X��
���8��BO�1)t	����y�<���z������9�C*J<{<�MwB$h�ƿ�#�x~~�mLϪن��/])Ѡ�e�%1�������|E����U6��	.�q){V̏����/1����@�Fr�/�YbY�<���(FY2*������X���X�V�?��Pۧ��=^ń�Z�K8"��3*
�e�Y�Ϫ��P����8-L���`{�]�ھw"y��o_A�Jؖ�Apt
�]J�*l��^[҄�޸�F���	���R�R
k����Cf�MT��_�U�q��<-16Yl����.ʽ�k�����T#_�BeOK��:@��~3�w��,��;;k'��e�ʓW�^.�4��&��H�N�>h���6w}����
bdJ�`^t��+�$��1��3ސ�7�w=�,�jƠ�)ԢƖ��R�2y}X0�<N	��';��7
Jg��F�d;Ys�l�ę��T�{�y��ZQ�=���m;���&Å,��9�",�9�Z�&�!ZI��b�~�Q� ��'L���8��n\d�d�L��%�^�L`PL̛�H�0��@%c}6�3�=ԓ�W�����r�_XB{��+t��Fh�F�6)j̱��	���?3Y�����ݝp8�A�m�5��+������W+�Oɹ��#d�@���b�X��n�&��X�0�����&��&{�z�m��|/8���W�E���pV#a���"�@�b���'����ՉdA�;������a��t�'2����̷';c�漡1r�&�#���%��,KI������[��K0}j��֡3��pA�<��ߴ�*liuO�Q�ň��$��0���ĪIP�p� O�����/zh�ER��x��Y9K�=�A �H�8���{�{6K����]X�T^l4�w{�p���{ݥ�J֎w �<�?�S�Ӄ�~FV����)�/��q0n�K�e
�v�
>�C��j�#b��_�����]%��oU�3�C�7�nb�c&���ׁ��K��!eh@��)���*���'����$!�O+\
B����S����G����p�<���'�s���aop��t���c��Ƅw�����a���I*9�����u�\��t��?�U�ڞO���g�C;����K�YM"��5_ ����́B�EC��v�Q(�d��J%(cX���n��5W�AZ��zvEl��YN���KC��cU8�c�lD�<װ��T[	��"ቮ�D.��!ID�<�50�r*�&ʰ�?j_�>UT�������=������L�%ܻt���Ǡ�K�Z	��i�A�4 g½������O�un2�Iu~4�`�epi]��Y�E.�l���V��G�� ;	�(��r�oj��a9�K��t*4q�N���n�5�xy�/��AH~%���X�c\A���>w��3�
Gf�K(��,�m�6��s��y9�����"��,_8�b^��0Bz)X�|������1%�1������!Yh����A:�!%��t�qm�C��-)��C`�.�v�+Mh
�����#6�u����������.fg�
�Y�������t��C�$����w�&��P��d&w�U��B�)����m�`�-����c�r��^Y�;��&��֨.'ʬ�!i3��mB�.�չ�afB8?wW��r��`%!O��k�f���2�ɺ�>�ʰ�Oݢ�z�^8����(%�2ߞ���l���Hq~>��(��=��[z_�8��V	Vb�8E ������K��GX�{�T�e�2抢���xwrPE)��v��D��!��Fּ���}��{(�bkך\���q>r��5:���*
@�>�5�#����~n���T ���Ɯ���VRG]�,.�J�5n7�IO{ﶞ]ѓ���;�
�(��f؅�s�_k�k�5�K�Ԟ�)����a����Ipf�����u.?/S�)���4Dy}�O`�ҤyLDzO��5��VB��lpi3�5��[�@e��֖ #�[�}�ޡh�w����EHy0������nW�Tc�t��)G�Ǵtx�	�,}��w�*ɗ��싣���D��ʭ�/[{���jD��@���v]��d���7�\J��O\���a顠l�>,���}K�(���aB�j[�#��T����U \��%#���a`p��@C�M�{I<�`˾��q�#`G@��q�l���"�˧�������jة,�ɛ��m��z
w��A��|���Ѳ^>�m��m��`U�3��� �ֈ@�
(��g�"�e`�O:��JP��dk�������`J9�J�6t=�״'y��(�y �fn�5]v��mua<E½;�2��U��k��`���yj���'�V�+����!�q��hhԏ8�}���l ���(��ٌ;z*�@*V�{���ښ/d�Y06	;��CtP�\��ϻ��r���X}�����i������zKl�С^ͩ�(�QNVA�i�=��o�[��2��7�����N\� ���r�3�vB����1��Ё��:f]���鏿~�;�E���H˃�a/�!z���k���, ��Ԑ�"�����KN����F���<X7l^
��{t(���.���9����`��x8�o����w}�2A��C��rds�L�<C�a��yS?{W#J��8�?���������4�,g�����M+�X`��=�����vJ[\_�)`�J�I9���u@���3�, U���_xO�������_JV�V�uNPsE�]s��^3|�{���U��K� �`�Te3��Ev(1{R�C��mΆT�W�+��L68�4��(MGq ?���!v$-���V�Ced�7��^+��7�f�'_b�v]�FmE�\�>�Z=j@!q�X=u��-�����K*��'�+#)<������b���G�0Q����(�#R�Z�^Ƅ��&=&�ם���c�.ϰ�� ��!�ˈ����sx��0�� ~�����N-�~|�p}�s
hK�.�=�6� �M�ʖ\��GS�EI >x	���OH�{�#�݆V�n���!�"�)u�@Q���`Y��'^)�3���9׵���1$���!�'�Q�	�8Ǭ�\�Ym��P��=d�r*�0��E��+V��XD�߀������|�p��1;ً�S�<��u�����8��}aX�G��5B���E2.z˪�8�Ž�F%��a?�!���.hO9^]�R,8��Hރg�钽�_�		���+Z�R"��O_:�>> �X������wRIq�a����	�!��9�z2�"8�|7[8=��d)=��E8�t�僣6���Óv��Z��S�-�9X�XT��p?du�6櫪':n�A�g1�Ŵ�����߱����; ����*��=�a��W{�7��`�1c��GaAd�qn"��=?����X�U�pYx�V���-���� ���LB�ᕃH%�{>������)D�^X_\	�;���6�[k�N{֕O3�o���"\=��ސ�UC�b%Y������I����W>c�p{{��1WJ�V���8mZ��O���j^`���Xa�*J6��#�f�5�qu�ŝ?���l+�}Za��Ï��S_S����69��5��.�	U�ݱ�P�;�$5�'ړK6Tψ�XZ��F~�:5�3�vL��Y���~ó�J7�˔s��2�K�W{	~C�X�U�tNo<+T���#W�U�̽5��@�2���~��"2���ۗ�U����Ü�ڵ��qEx�gw`պ�t.�T�Ђ�6Áli�}H�z�R��VMHb��$Ej��u�a��Z�>��1&\��>��jF�X�������X���V�k�.A)�/U	���U�� �.P)Tz�Ev(��݆^h�|�_Y����^5�q-Nu��,�,�2{�)���1.D�v:a�q�_H SZ�y���)���Suqϻ��7�[
j����ɿ��$���ى��%���Y�$��p�4	������b��N_r�Ŭ�+(�>t�w�q�w�^�e�:r�(���6�s���dLI�o5c�;����.˯b� ^#Pg�{yV�wM�X"bf�J�4�2r�:J�0Y��q�^�}�~�f�w /�-���d�(r��:�"� (DTBqk��cQI��͊��V�U�>�ul�JB0��n���L�I$O[=|�djr�(�*n
���P�V*�?'$�,ҨE��0l͛)oB=�|�A]��i�	������<�ޙ���������Ȃ����@29[�*�)��"�����{n�L<�9W�G3��H>Ɋ�BB�:�y���ހL/�u�p9VGg�@�-��H�-����bʟm(��ϙ�b��T8���/|1:�}��b�b:8n�`���B�5�	}
�x��f(�kő����y5��w"85�?���'�K?|�Jg(�hhd��#pF�#``��Jg�K6m�s8���X�k$����Bݎ��2�HM�Y+�󗷊fU���Z�����D���a/�PÙt��Lh�����.�Q�W���w'U2μ�g"�%�O7�L���e\��0��^e���M��M:�D�-�0�2��Pm1�O�F]�QS6;�m,]8���j�y Eϫ&�ǉ�L� �$������5�=�+9��+)���j岏u����9�O�u��Č$���eY���8��p���N�E[�:<���Fn ���r�����~�H!�����e8l�)?�	H��vHU,8�2v����N�AA�vZ~;8f���CD�:g!v��L�r���������E}f=0���kf���SV��V%���Ԕ�R����q=�8	Z��F�3�)�Ԁq��-�����1}]�����pv��
dZ�?f���h?i!ʓdmg8��A����{ܿ��6��)�eHW��'MK-�L"�r#v����/큷�\hl�`��f^� ��U��jF4T\�(Ep̌���U9.u·�
Է�af�9ɺ���Lw�o�n���V�E/[������Zb�����ɫ���&R�����-��}}D�8�7����$����?8��<qV��H�'��{Hq���ݶj���၎s{�����i�r��f��1�	��.����yd�s"�s�'k�����G�Wb�p�J�L�|�mUB���%�gƵ������3-3Y?��ګ�1J	8� �����^���U�\>�,��G�v�5P��m�<R��]f��p���{���<-۸f�s[��k�V�a��4�)>�9#���&�D�̥@����!�6��zckP �Lf<��Y�=�4/SE�7�h�S��#^���d�}�ְ���B�F5TJg����ꌩ���)���sQ����dׯ�|^>2�i�����p�K÷xZ��U�τ��0�V��!#�9����!Cb����Ma��A�W��8��֘��elw/���;��*L�<lҞ^��������)��nj�CL�Ecm��X����Yȓ�޷9����dB����	��a���Q��y�#f�k�#�S�Ɋ�/���|�����"���>ԧNj�Ψrl�jl�D��IN4�a���5�`��_)�>	eZN����hq���B������1y6tF��H�S�p���g.��t&'�7`���U����e����sj�z����[$�FxpZ5�.�9��s~�*L�U<J0暤zv,�!\�h������}�O� �#s-&MW�LM��[pϺ����^��P��?�*Q���G��_����i�3�y>9)���H�?m��.��8w����M'�U�"� �! *w�%6`CS�v�t=�8�:�Ņ�L�]y/��v-O0�Sy҆�nG'ƅnl�!�53s��5M�H?�P��� k#�o�>��5�{��p�:���<��Y�(K�G�%E>paӊ�bg^JN�1[y�"Xi*����f��s��MvP�g�!����@ɓ�1�L.�k�~�06�_��"���M�Q�����bT~VH��6���4'�BiYV`����aZ�o8�v��ІܳNcv��'#\�EJu�#��gټ�܃�T����<>�Ao*���@�%�)�꘎�@��`77V48������F�
K�~�(MU65ct����4��aJ�l���k�k�:_oQ�_�-�#�[ͪv�>�`�B��#�:�.���#����AP�0-�c����kp�*L �ڕ)�����1�7���a�#�������N�*�9SeÖH؇�d���P�
�V��|���`҆>B����C�TV�ՠӨ��/����,�yQ�05O,v��D�P�	q����M��F	��Dz���
���Z_�H����? 1��4��e;�9S���X�� WZk�	AL��a�7Lh��7�UYV������=~v��"�-���x�L�=1�X�A��ϡn�/�"o`�
=����K�d�(�#{��'�W���6��C
�5W��jY�����y����
cA�O��@�l`�n��+��VC�F^�$Mګ�5�[�R���a�$��q�E(�hvZ�p��1���򲛏��� 2��U�^M������@��������
�B�w�)�xj����~�x ����p�U���)0=i`��Z�|�A��-ڽV�;Rx�����k)GA΍�a�ϐa�]rb�P�~��,M�]BB���C?�W����]�k�K__@H�l���_��l~�5��k�A!l oAϩ���/�3m{�G�}���G�2ac�P�U�/��_˯ŊV�q��D�z�^�fA�v�6yȲ"{%1���N�����@��9Z�`�v%E1�9�!�;����f�g��oFE�w`�R���2�ÜV��e\��#�9@�a�f��?pH!�۷a�9�;��)c����;D�zZ����T�c�E�BQظ���G['R�<�r��4iA|����2�X�^���M���ܛ���/�hG�RN�,�$c[�ն�--R ��q>RJG
sa&���X�������L�W�:Q�����.du֑�<�*�)��uJ�ȿX��/9s2/���gL�쩏r�Bb�I����'�>��q��@1<�ceaH�8�3*� HX�}6QM2M���R�yI�_hN+ܰd/%�^Vؠ��[_n��-%��v�=ֿ��i�a���n{��WB�Y7y� ��tT5Lg��*�-�3k�8%�q��6{r���<,q���.�����C�_ɦw
�@%���N �G���4���XlxVHYEB     896     280��H�"`�$5�@��ݿ	��X�֌��V2cA�:>e4V���y��po��6��6���Y8�#�������ٜ,�������\����M���ʉ�pF�+��]Q�\��t���!N�I��)����1��VL~�Ű��A�P�4��Q��Es�����@ � �����Z߶z���]K�.��)<u���z�(�7n��q�8�H�B�aX�ɼ52[b-���� ��w��L�T�NY��p�2�p}���ؐHtԐ�*Ѐ
zHa��R9.�fy�*��*~���l�Z� �y��cH�:Dà����l(s,�A�XA�v��1h\)p���=	��{����E]M4�FcqP�F+�N3����T_��w���t�P6�s{��ꋜ���>c�;�l��Nz6���C�ls��l�' �!�iM
��\ے}��1g�ƛ��!eUN�0��st��E��%quڮ��K#�)�LC�=�}6-����o�'����/Ji���&\����'hڂ�w�e�����Y�v���ԇy'L����wq�yE���o>�=b�~�-����3���
�ݰZrt��Kh�����E{A��m���.m�0����8���*��<�G8�s�ݹh x7�}H�
�s