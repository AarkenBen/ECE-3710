XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������[t���Y�J?}�}G��[E�L�Z�6f����D��0�����7��V� �2�ҨsF��6�$�/��%�Do��F�&�7��U2'm��R&Y���r���Z��\��gOV�,>��DC��q.��
�SwB��6�of�O���Y��7ڀȳ�;�IKFeu��h�)���/�>pf�L	�,�/*G�_�e=j�I˱0&x�����"��!w�ה���ɀ+���E�a_G��3
���߹�t�Z���Uz�����B�(��dݡT��d��,[1&m�c�e�kt�Q�Ҁ��h_�)O���L���2=/<[�0�rR?�g)��F[ݪޛ^��O�|?衒��{Lb��X�����0���f��"c��:�jq���-�7��N?Yv�"�+l�Uo����}�u��Zu�ER�ȳ�қ��a�h����qr�Ue
N�Tζ���o<�濒��E��a[	1C�fٍ�"��6�Ӧ�d.��θ�p����l����(oC�Xn8��4���2}���"����U��Ҡ�����b��/D�-�oQI]24q����h�h��[1�����>C��vhf���£r�'�uν� �W��2�>�����61��I����#�M���nd�.8T<�M(��냗�h�������o0Ni�-���J��
�ǝ���;�j³L2*e�D�ԅ��!��?��wXj�d��tX����ϲ����oôdx'�X���e��s͇XlxVHYEB    fa00    2950���5M�S���p㕅�5��K�-�m��AG��WC+�!N:����}��	�?��}�[��(�ʆ<k�Ա����dNM���T�%J�,{�J,L�#CȔJ ���[�ѬŐ��2;5�Ю���ީ�����!��?vh
�5�A�{�a�;(��;|����kܣ����7���Ļ9rR�i����1�\������\�C�j ��k]�F �iU��6N!VW~�~%�p'�t5��Zj�	4Oԛ�5�畬� ;T|��þN��s,�Δ�r� ��Ct%��l9<��d}��L�#��ʷ��Ա�4��P�D�ܜ�j�l��^?d���/�\��kS�ⷱ�`< �c��������^J��r�|�Y�������Y�2m�?�r%C&�؆�܅0��`Bok:t[�#H �L�u���7V���F4#a
�r���|9�����]f����3��6��7��M�~�w���3dU��rGZ���]Q�^Ũr�l�pW[�/�������S�.�ļ����5y�(���t�	=�fd�RJ��r	i:��s�>:��]N8��[���ޥ�=P'd�wP��|��o�~P�iE�yHD����pX�X��H�\���N�>Ҽ@Uca�M>tꓷ7���w�������"�j\�vh���z쎣�+��O!y������{:u^	ָ$��Ɠ�
F�`ǵ�P��ȃ`"�\��fI~�Q�bB^.�bFO������v�I1alG����\�<�C�8=����>S���DiMU�ϢG�v�Y���n�ym����jI	���P�0���'���y]Mw]w�sun�^p׎.�y ��z�k����zC�,�%�����wy[��[�t]fmZ�f��A��{�O�+�n6�}��ڈ���n�2K��.�1jp5?E'R�k��v%���y�\����)ȡ�
;斢�|۸��`�R*� ��`sM�MM���͖iNit�2���o2�����*����U�t�$�jA�	�DBI7�ve�M��;n�u��O"�@���*��gn�����~�m�$��ÝԣZ�h!v���`�x�]m���-1� S�+�`��
��)?ARS[�KwB]rMF������lW��ddp6_��Y��wN�evBٹyI���԰Y����HK�B ���.рr��4M�{��YA�f�"{��r�Ƚ���7 �,����\�6]�c]�2�wp�S5Ro�^��4��F#����C��[�]V��T܄�0(�����Pz�>C4$����Ǜ�,��AO��E�h�;��n6?�M�=<�!{kW`rxE'58���M%��%�M���g
�E����p�bY���l<?1%<h���2񛌰���8�����A�]T���Y`��v��|=P��Z�M8�K�;�i�zft�郿���v]>�|�k���}q<��
��̈́���\���{f��������-xN��6�ng�׊e�z����ȋ)�f�g��oc�eOgmy�����NP?{��WsPr,_G4�s����y;���Z�,N���:I�t����fa2`W-��������m���@ɼQ���Q�ʫ��"y�ʓ�?b��i.�?#��x]E�𧞥��F�tǄ�֜�8��A�<����L�U��ʥ���_�����U^��Jc-#'�0,J�P�o��a�	e�2+�)��Z[���ŔO�c�TJ������+y(.�M�4���aY��(Q�29+0�D��1��NJ�N*��BK7ÞbG�8��#nr�uzΫj�_�����M��T`�6�c���K;\&$�VL������c��|X7�I��+�>�5�sj�	��H��7�hm%�'2]G�PLv��6?���*�0L�GV��vY��i$l�>�q�>m�\��I���1�����#T%|J�s�^�_���Q��4j	�Jc>��k��Źw���®�.)�b:�+�t���� 0�hT�ɿ1;?/��\�<��1��#_s"�)lf�m'��7ƄN����ɕt6v7(������p@�&�Qrƶ����K���A�lJ���9"Ì9m@�+�Vyg7g|�#��L*�ߟB�6F��8��0�[:z{��h	���mPpN��Uq:Εo�ȑ.W��ߣ���f�>���x�O�n���;D쎅��fDY�l��H��B����`%D�������W'�V�Unh�A�N����F��RU���j��n��`n
�����|���LH�t��q�V����{��M�5:�ek0�10˹����|�i���N;��O8�|b(�'�u*��ͶYL�(�
�wS9��_ѐ�8�e�������:͎{����ò�/�жm�2�jdl~�;�R���$Þ9��/JP��.����@g��ծ��j��܏	��9p>L�<�\bwV++���Zˡ8�l�y�e�A�Uf:ci#*9��#c��&Ü�g����"���I����"��~��m�S��Ա�˔um
��u���a�a37C)NCp���X�0pگ�0̟�˒=�x�</2��6�N�;A_S����n�m��zH�1��<@������\Ld����p,��>�s#w�%)
��ݓ��K����=	�ʈj��3��f��lABn5FF���u)�w�j
N[\i���v�z����n�.���8�9��&2l��
��qTሯ������6T��G��R�g����r�dDqތ��<��~X�ǧ#�i#��	����p��_�'��hIC,�"R���h��Uɞ�wB�iAU��p���Կ~(��/[B���dmr5��S���ww-0�(őc`��Ho�g?��T����7�=^懸AgCoG�SkR�悸���L?O��'���<��ד�T��S,'`���3���6���17���g��đ�|����U��P���	�I���_3 :��y`�Lg��N��`³���\�E�)�D�쒰�@��(��R�C�D,u����۷x�p%�Ф�I��:G�i3:�ܲ*w�k���}��@��{I�g��^X��jt�4vX��mCX��&����[��t8d�P�A��]�~h0y� 0۽��k١]��D�!�� Pp-&0�-l_R��=���P�{U�D���\����o�(,V"�-��gZ�^O������RG�G���t�+(�,\��N~�M�>�#x0���}�.��ɜ̺YΓ7S��4[�O=�IJ��?�5C��an%�W��4�U[\�+l�w�� ��q�z��Y���|f�$���@�Q�3����p�b%Kqq%qC����j��xo��3��!ۥՔ�^A:g�MH�Bҥ��f� v�yۖ���g�s/��Z��B�0���p�!�����a�
���F5Ĉ�rx��c���?� `V4�]�0_Gi��Q36X�Ԕ�t-�|b/�r�H���b�?9�����f�@:�����b�����q~�mV����`�m�s9{�W2qm����D�,�����
��k��t߾�����Ѡ	�І�0��\��5F�|{k#g �I9/+��ڂ?��n�,N�,!�E}�k�g[�l�A- PJ�T��bǞU�¡�tU�^3 �2sCy�d!�� �kZe_у�x-D�S��Xh��"j�#�brA�vZ�(�q�EqJ��vRҵ榛j��9�Zmڑm5�-nS�RF2Vёo7iq2k��;�B+tm�;�ͺ&�ir t5D4+����\2�u�w��v��=�
�d^���t�c��tŅ��82A�&J���&$y�#�We���e��o����b��KY���R[��N�>N��э��^�G'��%4
�W��*8>[�ᢧ���Vfے1ȡ��#�K"�pBnԑٔJ���LZ�W�h_��1��]<e������GS�i�{�i��8�%��3�/c�i���Np�Y��~����0o=����)�<��^��@���,� �����r��@˔S:��F��3u�� ���g	��$f�+�Q(�y�Q����"^�u��8H��k�+Ǣ�h�R�F$6���{ �0��W_��Ss��p[�����UԭK��Y�8��T�@�D������H��i�_���k�B��������V(���m]kW���.�p�������S�{׊~=���{�ڻ��gt��p��En�̵�KBl�;k���|�C8��l�/8A�oR	�Y}˄�r�x1-�³[Q�L�3�uܲr�����
��R����UjacVڔ�m��0�wܕP��۳=?��Z*��]���CMs��0�&�׃����"��)1�"
�eec�����Yv.l|sk��'ۅ:��W�����Lz����5$Ę�^q7��Ϙ-�գ�d�^�uФDh�<���G�cU�O�=}�qk�sˤ�2.�t3��T�'u��A�@Z[dA&�g��n�D�b���&'�Ս.Cr�x�qo�;G�!3RGY��hD����f�3t����T�b#̾��q��̜I�8#>�T[T܀�p��V�l��V�nk>��eB���ڐ���Bk>2�#�9E�A[;�v��;3�ZEE�Z����<A����i�o𡙟V�8X�FPӬ��D�˞}FV�T��;#m���N�L����6`�� ���B��o�D��n	���R�O�	Ch�����o�f���"���B����Ec(�n���2�	��G�T�2t��{���%����D�Y�؆˾7�Cm��]�k���P0��uN����]8����E�ൎ��y�%K�h3E��5��H�%�N�(J�TN
�3�i�p|����[h/�_�^}�XQ�O�B���w{(:+DƎ��i�Ej��A�۫::s�.�;L�D���e����n0Ɛ��� �e����菕�M����N}?(&����$�͂k�X��Ed�k�<s�ݶ���R��e�)��a��z��.N�@�3�x8ۨ/�[��LL����fX:n�lhL5�w'"�C�!��J��tj�������oiZ�9eh> �n�ͽ"w�c��i�r*�����Mb�>A��QpQ�{���xب�us>6\>RX�n3��2�M4�������gtn��8���*s�aW���_�nI��΂�]��������Qj�<#1����Cp�(��I�n1��-b����1���&UG�ዏB��+�S���G��\����,&!Z_��{.�5LSwt�LK=3�Wm�|�˛������p�ILl�������R�ޅ����@�$\Տ���Q#�-��EL�?n��>^.�ɂ	Y��cڌ&�I����-YCֵcջ�M�YFy�d�Y��:'9߅w�s#1�LF	\4T�q��_�S������`E���|���Iw�G`�4� @���"���4�B��i�A'><��BV3�+:�E!�����Ijz4د�5O��O�a�x$��[$�Q��F�=/��Y��e_���<$��&��$��+��уWV
Z�"��Pљ�;mdF�g;� ��^�T�##���L�֒�O�d:���d��q��\�����'�֢&(��|;�_!�I��Ź�7k�Y����<��`
��:������A=稏�ϱcv��$�g��X�����|����=Yn^��f[=���ƃ��H Nx9����o�4E�׆��B����;�4_7�L�'�QN''s::���	�(n�����RE�Э �{}"ņ�)�X��Gŧ;G���l�FΝ�*�a�(7:��4��]/WmK�
��*tc.�vX���\�W�@�(�&�~��q��LD���s!�W�Q��@����Xt#���݉W.��<`9�P/?��������,�V��P��R�z�l.+����J������Q@hv���#��@�G P´ �wυa U�6Z,�E��4j*A��o���e�X�a���V����Y� W0����"�?�E�fV���b�����`�D�U)j˳U�����b V�JHV�(�L��9����8�$��b���'�h>v}>G
��fk��l���������Ag^���6�h�����2Ү�!k�ߟ����>�ByUc-���%冀>�.�-�e�y{zV�ay۩\��	n����K||��!j ^Oƾ~1�H\�[� �R�*k�CgcZ�]m���I���4v�a&�/��tlp����y�1�N6<p QW��pw$%���ӝ����$
��-�/G����	�	����e����I�J=�����NE~�Y����Ⱥ�Y�@Е�^	<T~�g�)��[*�V"%M�Q����ê��@�j��g�-V�\�ᨸ��ՠ����l�J���=��<#v���������Ї-��m�2�@U�6}<#�7�M����Qu� �/�����Y\0�R�	i��N��,�	%˙�'���w���I����%_�o�������A}��c�d���_>a�W�oPذ2	��>�$��IŇ�eې
tlܠ�/	�*ԗ��4��K0�R�n��Eլ��=P�Ai���S���	̳z�*�CsY��CΚ��$�+W̭�DU֟^5�Ǣ�-�����"��O͠�������}�5�hͱ���A�/f�|�c�2�:��gv�f�L/��`aR�L�od����z�SleS&mVy��E�BRt���\<Fw-8{��N�:j���V$�D�T6/(�W
/G�E� {e{�΋4���3s~�`�%5�8V�+ǻM�&�`1� �%+J?�>�����=q8ۙ��=E,�-�FP��H�'��?�2'K��E�U�s/Et���`��y`�H�bfç+>wa4n�ӝ�1{Թ�M�K"�	��3�9�Q�:5��}� ��e�E���}��U��3�5g=��6�/���g�l�jI�#;F��fK
/꽘�[�X�����#����#��C��m�Q���Qg�p�����\"� �3s2^��1o;�i�ڀ-`)��|��Dh�����"�0�C��o*@��d$0�#%y�
�&۫��j������ v8T���Ы2~��R1��~��ǼfE����!��wN�,����nA��� ��I����9����D�E+�p͟]�Mw[�a��rx9x�8|�l��r���-�+��ophme�5�\�a{x<��� �a:�N�,���E�OL��V���5�F�2�����aY�w�Cx�G���s��& �R<�hߨ1Q�R7���S��U3�C�.r�ӑ(���q�_!�f�R�����\�����t����n��I�t�=����Ҋ����+�܍�kD�����<aYER�ۇx��7���K���=��}#k���oHbAڽy�q䇹x��bȊ���v����Tѷ�
I����J��������������2/��+Ƴ��v3���`+�賠�)��Km��hDx��P�/CI��Wcy��u����ZS$��1��}Z@��U\�n!А#�Z����e��1_�=�/�&��&���?Lw.�-B$��S0I 4ٜ��WS�e�4��DAp*iU������O,hn�ې���'�!(mOg弦f��l�?��a��$�۞ ���#p���?+��"�]�9-@�$�cv1	�e����Q�b�ļ�y,w).'��h�;Qv�Z8*6OVd8��O��a�/k��DʂpY{1[�SЮ}i����++j� 4�A~P�&��[��2����*u��w�ldr9�9%��"�x�&�Nl�q���qh5R
XĊ;�Y��U���� �m�4��k�$/����=f�|���'���;+��y1�_	p+�q,��4M��p��N�}r�Wd	;���aj���q�f������������`�  �o��<� �G_�4��oye�)P�Cb���f�h�G~g��Kw���vm�5(��i�'�2��A6�^&r1>^nV�@������)y+�Ƌ�������.d�k���u})��g� ���2C�ד���b�.���|9�L��u*��@��J�Y�p�NŇ�2u����1st��
 G}	��㓉�nx�K���a��V�g��YRݡYw�����R���쮉!#���q���P��R�x�ǼF����ٝ��elk��F���7�3<��9sre"�zn�yȪ����7������+���w���.
SZ��8����i���ӆ����D����2򔓰?hԛR��#aYؓOh��ez�2ؾ5f��*k�"���?��&X �8ړ�W�(O@������U�,�ѡg��{ Ȩ���p"?+�¶�^�b�m��ܾʦ%kD���7o�S��A���t��#=۩eK���������w�0��?�j��D��@���Y��*V�����N�o�a�������!!/��m����c$FJкzQ�����<����F�~��t����8�S+�DT�u֍�Q'�gb�L���A�_�3fF�J����j���SuL����A0������*ϟ!�!��qг�)��b1�%�y*tM"��n'Q�pA��4]^u�
]�H�<��=��W���QŅA�GR��|���Ʀ!��_�����+���@�H�t\��\�c�Qmr4�Uu��-s�+aN�Ch����羫E/l�WY-�O�~㑯	��E2����ލ�t�n���s�gY�nK硈���I|P@g�T����c*�.XVd���Qu��r�U��+�&�RS�k��e����LƔ-������������� Z`w�dd�ͮ��l���刴�Y�&�W��ɀ��~8�#��ք��i�[e<��&���Sw�����D��$�aHuo�d\짂�(�#�Z��GN�P;�\��,-�.
�����mp�q�MEi)�/mO%���My!��RF�C��
�^[ɜa�y��f�5���b{.���~�u�E{+�2�����/_�F|sM��ޕ�����b/~��i� êkqb�m����U{/�l4F�$�z"������V����)�B�9c&seB_N�����I+�z���|ڴ�#��(5�����C����q*�#,.<���>s�/��>F\D���G�Yӥ�k�^��4Y�(�`0P\���h~1׏�o�)duפ'F��=ԏ�
߹�S�p�%��ۣ����D���4}Ɗ��t �OH�E�fQQ���~�uo�f�RQMv�����[�����^l�J���J��n��w�-1�C��Fc�B�d�'��!�4*��I��N�<s=-i^,z�@0��M��1�p%��5g�LV��o�a�Y��(;.Z���B�A�[rP��8�H�dL�_B��|z�u��GB	�:,�wV*l�B��]o�����E�l/�Ư�j��7Y" aAxCo�	`n_�����=��9�N����T����^B�9\4�����pǇjt�Q�QnOwH������A�a�}�H��B$}����n�fq���&r�+�`jp��ذ�T?;�(ƺ����jEӰ��𼋯g����)i
U�� �ׯ�Z��]�^��/����DQ2w��d0�#������.^V0,:q�D�����a'K&�Z��[�a}ռX��<��]�A�g1��6%�o
&���q�IN�s����z���ԅ���ك8�O3��i����� ��'�V8CD�pҰ������v�'	0��ذϻ���a�s�}�TP��_�����-�<�N8X�Dp��+xD���ۺz�{�	��"P~*��^��4O��z@­�I����E�Y��4^��Ow,ABg����1!��L��P��8IL�V�~�ѱ�&��l��UZ���>g��sK^Y�M���6��R��������"/���֊�1�p�� ���b��\o��O���~�"�{7���E��2zW�M��	���nH�GVL0�.,b]D�7�&�T�D6�R�(Χ����z�c�~������S�L�I=����9�5���.�'��@l��	ǂDX�~���m} #%���1 /��[ �_Y��-��lT���Θ���j��u��@)ll�+�?�����آIH�XW��l%����]���Ǆd���~�YQ�mw^c@'4i�}��H�{Ķl k����QB��B���:�O�4�7q�!zz���r�F���B���Y�#���h��~����=�gݝؐ|@� ��ӥ�Yz�FqI":S`f�͗D���f�K"�>Z�_�U�&��:�P������ �1K��d"
`Y�%������
����#�ˮ�ܬ�4�q��ʚ�����Sk�}����8gc�������@�ڊ�Y�w)���`a�d·����JA�:�Q(�_	%عI-5��+z��aCPX��7��7�m�X'��v{>�XlxVHYEB    fa00    1e30�xT��I��@������7|����`b�v.,��s�g���g�����f#����5ڧV轻���[�#pD�<]�6��`%���<��T ew�\�����6 Ô:O��}V���1�qE:��(�mg�A)��m����TO:%�e��h�^x[�ň<w�H����@<�жF 0z��u�/��9r^7@�<�i,�!���nP�{;��P,QzR־hx���kR+��0=� RUK���_rp�R&\c�D��?Cdo�m5�L,�}_�ŦJ����\\�A�]���_����_�9�p���$��>t@���^���A$=H�W�1�Y<�*[Z5��/����m�MMi&���p�H�eˀ-�S$Y��+J`�������@�/D0�4w%��d>������D���讝�]�<J�ŉ��T#2��wVy�b>������ѡ��6�N�P#�����'7�L�������$�H�p؅��S��a�Ч�G@��]���
I쎹�bI�X��܆�b�eJ�oßT�)OI1E�m(�_@�p�01���+gܩU��i��u���ē_�I^�	���iBI�,�!!�l�@1�;5ɩ���C�"�jb�|٩���^�G��n���9�����H�fK/&��}s�����������*��Rz�1��6��d�t4o�����V��G�D�V�Ѿd^�8���'Sft��xf�*�C���{�Kp/Ͼ�o�'?�a\�m�fp�b�%g[���s�'�|i
�{�n�TGe3�
�>p]��9�����ʿ��[���]V����R����Nrs��&��c���j������6��(�p����D*��S���#�Q^����g�3tU��*���4�0lE϶�PK�����I�+Lv��ߟ�.�%h���EpZ��.L��[{笤�MI:���F'���Btd,�S�7�T2�Fб/X�:%;�J�؀<jRt�mCBY�ZiW)fXɒ�L����U�,ᬝk|�'�ѭ&8�U�@����A��E� �u��2U�h��;[g�l���g
>t��$���b�u�7@B��`k��)�GAE�~T�G�}�T)6�5�ٖ���q�8B���H�aq���a�Z���:��m� ���yM�Y��u��
�Db8D	(�­ ��\���լ�v�0 ��r>qСh����y�
N7�+ �S�N	_L�*'g�	��qF��8�о�� ��R$�-M[i-	L֔�R�"裵�Qf�B�ת�H"��|@�^k��m�8��!��ȵ�:�?�d2d�i�^�1��ۯ(�="��ʐ�h����heߤ�PԮ�Z��#���`/6�1?��Vc�R��Cj�1l�G��w��--N���:]*=?t(�KB�,���)��z⁗����Tۅ�Qy���%{AOX>%I�?_��T���z�l�>���9"b�w0� ��t��Uxe��Tޫ�r:*ٸ�e["�=�$| �MC��_� ��ا^6����7`���X�Z7���d���4��] �c� ��Yؗ}`Wx��"�>/�E:<���mYK���D������Ӫ���u&�o���J|W?�<���3:��ƇH|ѱ|{S�ɱ�L���ME�\�^�1)����b�����6���#�����+L�գ�5��8su��?#JQg�6��7��&��O?�#�3S^�YT����m͢�SR����CW$�G��
�į��IY�8��
K��ǌ*�Hq}�4��<y����"�y�~��:���ZVG�+jD,�D��ǌ�)x�*����@�>q

�-�8�yĄ��;{��q)�0e�f������Ѭa��)�U	-{�Nx�]��J�u���6�y૒���������,���z�T������D;V��X�޹�?�F��c$JDtUE���S�6)@!%���?���0
N�B?>��;���m\��x�kr��<.
��o�E��<��R���(J��m�Ы�:Z��.�ݔ>"Ȋu�_���^���m�8��8r�J�H��<�˰���@7����,���lJl�fɵ���d/^UYm�;��G���2|~+l�}�K���P��3fOkb�����i�ys�UˆM���بo���m=�vm����p�u0��������6����ײ�Buzd�3f��%*V5B4�ƨ��JJ,�A��)�D\�N%�T���5��V7�M������Ltu?�@`����Ci+*ow[w;n���k^�"/�@/"ow]��n�j%}�����nT�T�T6�산�3��k�/��+];�鞒�-���͙kRhﬥ?�x㳷����܍ȩP�3��CE�������7�b�)aČ�F��f�[ފ=ӫ��p1�=O��n���=T�PH��Ikt��2�7��x1��Ul }(�G��HO����?�@�#��)��g؟%�;�jq��e�\�
��b�c�tKΒѣ�p*�-A��9u�#�Mb��7SAy�ᛒ��"b��s�H���M"�W+���=���I����4t��D��9�̒#)|��#2%�2�0���q!�*ۅ�T/�)T7�c/#�����tMx/�◌��i������ߣ������2M���vE�YryI��M�4	02���4�YaP�B	���8�'��T})�|\� �n�q&���Ћ�V]�����<�:�y/\�Dix�67��DO�mV$f^��T3$<����|��|��=����>��8��V�%JM�7�ќ�o�T!�bR�bw���~Bnn�S��Zg�����:O�\��R�m���)P:0re7�y�8CĭV���C0�����Y���|d�2�f�3�A1���aY=�X��6j��V�่l��n��[^w�^�E�DU����-G�D�?{%�p�u��g_t g�<�Z�hj��Uoԟ����Rj��H�T�}v�ݞ�}N��W�;���P��k�c`�f��=6��8�ym4�.����������x�>�Pr?�F|�Đ�8���q���wAGh�s�U����|�,��@'B-?���d��g�Zu&��GP�:["�':�<j�ո���zmN�}:�=����c\�ܴNxα���3�h$�;h�7�V �V�>�yn ��|!��M�P�CѪ>�u?Si�o�������x�
�B��n��r����p{&��X�Q�,�->��8G��34G5U|i:w�Ȩ������{z ��=�(�װ���;����9<��ؖE6HġMd�`zm�c����M�s��Ҵ;n�K�F�B8R�_�!���P~:p���%AZ�c�Z�W-��JZh8�:F�����0��X�9����ϊ�佭r�^J�H#��6T���zz֯��X��e�R"	c����\�j��]�&�	>��5Mғ�l�/�Rʑ��e>���t�MCϠ>��e����`+��p�S8E���{V�Q�����Ǘ/��t��'�I���!>)���5���(T��Ĵ����r�j��bǶ������P��D]1���)*ձD[Q�m���h�r)��"-.�]zZ�hS]�e�,(?iH���p]�GO��g�X���:��h�ꏣH2|5Ze?ȩ�w�7V���5�c�xKWo|	��Oox#�i���{�ߪ&�ڝ9.��ZA��(�-���S\P ����kp6�F~�x~@�1����sm1J�%�0� ����[e�;&��>��[��v d�j�����ƺ�gvd"�����HK˪ efa]�1h2�8��v��ǩC�������"�X��?�DK��8)y�1j�"p0H<��@�'�_EX��܆|����2p���J!$
5�G��[�Q���5�T++���>Zᷦ����o�N ��ڣ'�v3d�?7�`�@�� ����p�E��w��U^�jY��ރfZ�u�J�Cyn#���^P"FwQ����S�L�#�>y�0��g�h�:N�U�I�*i|j����$��r��y��^C8����U̳#�
|�fښ�R�n9?T��H(�cM$����.V�}k��$���_�����H@'c�ŨB�\�J���YHa�ʜ���3{w��l4f�V�U6�GO���3�3�7/�:��z���߼��1��]-���.�k��eJe�W,OP��s�zF`�o��Ne��oM�l�q}Ո�. �C�Ҙb2D����w��U�כ�)�S\dX�l֏�B�\p&I��}t��b��X�O\d�w����6�&��P��op������:T>�'�6�n`����X9X�3C�~��2ZE�i��N�����H_�G��e����xV(O��@�x���>3�?JzG��g���\b��:��zFK��&�t�	����RU��8�;O}�̀���*�"��YJG7��{���Wg8��w�1���'k]O~\���� <Q��Ĩ=<�0�7�G(����O��qJ���6�E��!!W�>Q�WQ�]1�_����z]#W��#�Vm��C{�L��R����
ϳ��RtZ�"��?�/�^P�*��]t����To#���ET��F�Uc�J|r�ݕF�~�Zg�~
���q�ۏ`Qb2�D�iu�;A��E�5��N�~��9���CI�AR�pOSZ�8cW6��]�k�/lU@���7����@�u�Sӌ:T�|�$���	�Gx	�� k�����x���pa�I����﷨2���q\V>c���R�Zල*-���#0�Ͽ���z����1��jո7w7ی'EK��R	�(^�$x�⸟~k�Hاnw�o�+ؐ�t��E��K̙�tN@/b(�3Av�\���U���jk�C�(��%x&��/?Z������Y�jp�x�:�D�0�ǝ�"�a�W����(�	��H�˅��ӝ"�C��O���x�>��h�.���%��;^�W��
������I����C�-��1]t;���z<���A��C_<�.�\�j��z�3X;S�������Kي�M+���2��ği����}d�9���Tޤ����I�y�܀�UƓF�*�\K�a5�N=�<�&!�#���c��Ј�'�xf۸�ᜓUz�L ��(�̼Q����knF-K�}	i��j�VԌ0�f6}6�S�)jݗ���LiIr������)��1�ڻ�ԫ[��G������*;��kKj���~��1�`[����`���I'h���$�X�E I�dC���g+�XA\ɳ���B����O��s�P���eԴ䍛9��`4��q36�K�Fo�:q�@d�E�&�o��A�78t�����*�	[]L|n�r���د���s�b�v���LBG��[E�6|��Q��*g������C:�����,��!�Ҭ��{��;єf�S�O�����(�7M{��Εmn�=(U�D\���tUai���ۗ{�;Ć�#:8	ďV@����)/��9~-��t_��S�L��^D�Gˍ��!����(��3��٭���\f�Z:y�ɐ�\�>g��d��C��)�%�-�z?�mD�|�t�t��S��.�}��NO݇�{F�j�I���C��|����J
^��3�K!㛭n����,��q(J�9����TK]jɧ��[S�M0�c�)%x�h{^{?Kz��S�_��I]e��������+�#����/��-��eV�QU~�d�	ぺ���F0)b/�$����j���}w��xq����56xql�s�fuBS1��&%��	��z���X�g��/�!5��ֱU��Ώ�W�c{��`2��K;�����c�y+qo��8�(^I�y�����f+n"aA��EPQ�r�52�㸵/~��/
��/v�$-:��?�ݽ,'&�P�/A��^?��Wҏ�A����0��8�?n�����rٝ�a��=G�[� �y����XS�N}����/��/wPO$��@�b3fb�Ą���/:��r��Z'M��'#k1�ˍ�ro�/�jF�Y����WF�yXhn��e�� �
��˝�h�+��q�;��eB���:S���v�W��ƭ���üX8)���
���3����%����5��X��;KMBPE�_�!�&���	��mF$��� �a@]�L����v�i0O�`�ki�Gmj$V��L@>&-����#�QF����eH�]�Ν���S�H���w�)5.�hMW	o����=�_W^������޾d�"��S2�~w�B�
��pV����wDz�0k�>����<�շ�;6�o�kA������	Č4~�C�Xb*p��b�~�QR�lSV��������W����M�z�˖���p	��U!����U|;/kb��-=�e�'d��Y����W��K�`�:�gWXּW���ͻ�?��o)i
�z�lus����j'd�
ҏJG�E�B(�����%.r�kM��Q��/��ڜ{�Y��R�<I��?�*',��E�@�w]Z_Sk�S���5�I�e�&�J�hv�0��v�r%u#|�����-��(��O��z�Ƕ���3Ӥ�9@[SI0���d��v��k|��غ��j�\�{�{�oGo��)�/�r�
<�S/��sLqh��D�,�^"�rI��T���t���n)y��a��{UrSX�4����T�����J�w	��b�H�0R�!��:��(�
� ���&�����Z���!�ʁ$m�3�B��n�M�Ө�w.3�S��e{�R�إ�W���{j�ug�8h��X.W�O�;g?�(��P馏��<+C'����$�~i�������ܧF!�&��t�k�9�J}�$�֢�)���;j^��R��#���_�<���áZ�4A��X����:�v�贾 ��B!�nï��ֶ��'��ob�΍R�z�Y��z4�N��`�}7�Ɠ��xf~&\1+Y>��E%�;ͭ�#Aj��?�8=�i3cO��~�Kuk��$�m��3�K]a�g��	%�kd����R�3��A���&�"��ʖ�%u�*LW�n���̬"������J=�.���2Q\����5M��/ok�@?����#E)��. ��ϲZ�:&���2���7�:�<I���|��Q7�t�x/Z铛Qa�PI��">��r?���K��u����ћm�� ���Ds��hm��7�[f%F2[�!jfo��o��A=ߏ�z>W�Q��)�'ak΀wy���*�G�n��^Z�'�|��2-�0�����;7n��F���kdL|�if{Й���r�9d��ѳ��@���T������*��nT��H�ˆ��S�^��E�.B:�@�D�:��=t�Y�����|5�Oq�xEN�e����J���"�׷L|�p���r�H�\.���$��K����>��QFO��e������z��	�0�=t���=%>���W�X<��v��S�,�AՂqg�/�\k�Uj�5�7�,��&[1��w���V�I�S�� ����C6�a��B�-�XQaI�f��E�ez<L�c�6��{����^{����Q6v���V0q��y�h���bp�)���L"8��鼭wp�c���*�g�/q���O�-x���&P�+w�Jv����uf�˛%|�o/XlxVHYEB    fa00    1d20
	c�_@Q~勮�Fʿ>��A
Zœ���Yx%3�(��aXw������#j[ÿ�G�<�v���OO����*�|)��:ڰȱ�I%Z���%h!����!���U�����$p�4���?����UtNsk�{VK�F�΋����������D�r�qW��8��d���e٫�K����:���O�H��W�����;u���[ϱ�pk�j`��6�;t�!
Pm�K6��S�SK����%$���ɲ��{B9��=�c:|k�dV�B�A�6.g��kt��L3OH�@�D�%ȅ
�K5:��|O�ɩ���(�O�W��|7�� ��)uPq�T�mǲ�O�u�J�GT߬vꥋgQ�������s�e��t�-O7�G�����g��9~٥�a���Č�G��ݳLZ�k�R��� ;7>%v��K�g�SqI�tG�w�zhNQp_�-���|�����j��.SA(j�H�w�Gp��[,���l	Jdr��V��[L�7��25R\/ʾ�?@r+f9�^��Z��@o�aR�fӈ��djc��3�TW?�G\tN���'�)<#P,c^�e���HM���c�����6N6�h�"Tݚo�8U���9ԫ�^}��45Q��=ID�+�4��W�*���(x���S�ҿA|yK��[�R����7	�[^cB#s̗p���)� i;ᕞY�1Tǵ�H	NA��H�|i��Jx?M������q��:b�CHy���:K��ĐAy3����%nϡ�b-y��4ߞ����[��˱Ydml|))�&�o��A�o���W�Z�po-0 �Y��j�As�����F��������*4U��9��`A֣��vDq5%�*@��,-�#�k^YD�����������;��R�"(U�<	�{Q(��x˿���T$�~t�i���e��x, q�<[`W���Ƌ�F�T�+�ܲ�9B�WfG>���<�q-2���o��2׏�U��Y�M;5�,��Z�/&x�cZ��Ϗ  ���ɷ>Y��m%�໾ ���A�o|����y
2ۅE��#Yȧ�5��aº0˒�Y���xd�@0
����s����!��H?j��革�wV�@Arܿ+eN.7��|L=�Kr���%>m�:����}�a���+L�cm���9[{�k�g*�]ov��3cCq	�L�Z���i���*�Q��1U�0N��J���΋�3<���L����5�sX�F��(!D���&Ç����w���_1��䉶y,�Z��ip=��1��DVv�����zA�Hثu�
b�z�-Fj�Nʃ��(�z���ɘ�<t<��i>�.�'"��du�(�\.���;������b�"5
��){�o���n*K�~}���FBu2	�<X�<� �o���Bl3 �ۧj�G����vED_�8;�#�c2��Q�<�ȿWԣ�Y�<�̥��c֡쀮��~j�*F��>J?/c�k�U�,������;�Y3͝��1�D�z
r�`�8���'�k���c
2���'hS�Zi�Bӥ� �8�;C_k��k�ˏw&$�� ��ࢨN��k�n�cUMS2$��v�~ �
�]E�[�2��杫�U�7Ɉ�'�O�P�z��i�1���ZGC	>��XE����hy�ߑ-<�Go�?`p�]�~u�[Ef�è8�ݝ��ƙ�μ�;p�GlMFTn/uԧ�gM/��p�h��s��,�5�s�p3PR�
��@�g/ȷ9��D~�T([u(�A���?1�_��i��Nh�ǃ�������泰n:hY�%'��`	,����2H�um2K�H0Gdݦ#o�Z9:�bq�H���������`���{�=��˽��g��i�����:�������+�;��1�����M�E����~q�5�1��'��O��D4�RJ��%e6+��A��Hك��83n��>�pZ�J5����	k�O�'�����<��:(˧���Ev�^�'�^$�2d5�po��+ޗF]`�?G����O|�܁ې3	��êl �	1޿l`�Y�X:�^�n��D��e�����7RgP��7l8��:���Y��Wc!�~t�b�)��44�ɇ� Y��G��C�'C�vIG����?��7��i��K݁�i�S��]a H4�m��q�]���W������X�9B�H��Q��IpaN�ƂU�b�"�����r�@7f!BQ��)����z-Z����#��45����И� �����+2��ŧ�76��d=YPU�Cj�0g��8X�E '�[�!X���4����OU��?e���{)�������
6?/�>��A֪�\qG;�7�z���WIY��n��Te���zmK _�=E��� C��f>[Wp����R�����Tx���7�.���l�u��hLa���w��~�^4g��ƅ�[m�[�,b�cu+2�}��Ig� B~��#����Y�Ą6\A=,��_F�jdN^{����NG�[2;֫n��1���3a�����/*�P=��J$0U:�s�cQ0�8�i�:�R�����TBiӍ3-��$I�_��݃T�K+ѣw�x�{	G���xJ�,wISx8�y7�|mDN�|#r����ƛ�6�s�F.U�kR�L����G��zMO0�!Ca��6h ��~�V�G0���x֚�X�=��m��N}$����0^H�}���\��"2��]�D�$ތ�W��! o�OH:���N�I��k��kft�����I�d B���B0u�#V��ᚯ�~
+,�(c~�ű�U��gWEmԅ�<���iϪ9�t1; ����؅6?:�w'�0w&~(m"a2��
��Р�Z;͗����U|�S���f�R|�򑙘h�C��`�D[� Q��$��vDU���?k�M
TE^�7,B���U5V,i��V� #�Y�A���q���F )ŷ��ue����_��i�!n�ٙ��=��$��3�~��k�㉷�mQ�<����W��&s#���Zn�z�HL�Ŏ�be.�[��0�
,ﭺ��4��,�3N-o��M�h_�M+'�����?����<ww��4�]�v�5��{�Q���d���q,#J��,��|�Qb#իk/��YRl��\��+��1$��|��?�r�T�!V������
�M��O�z����ٌ����V�i�Pr���������(�銄2.5�7Z�ږ������E77S��87�V�;�ء'��n<���fX*���>?E"x><A?�#۩ �bQ�����n�M7��(5�NE��Ju:5��`�%�9 �ěKi��¿~A��D��ķK�:[�w��ț��LV�	�Eڍ�^�������e��kK�Q�7�`Q��27PCZ�Ӯ�Y��Y��޹z�s��97�q+蕈C�
=�-.�5����k,���$�]��7_w���k����2�dfu1�lZ_�9ANh@�XA]`��4�W��u&q��g�s8����=)�2��1��G	�|�>����D�}j>@,J��B��2�1.۞���6�]��>rt�����j�K�~\L��:�i���w&7�ѹ���Am*�u @o��4�$�Or��I����@���?�MX�"�&�қ�jv��A���@�9c��G�GF�s�P�ǿ�O����p����*F�Ñ��ܑ�z��l������:lB������(����޹
5���o��J�f��X[^ kG'G��R�Tc�5��]��ӑ�����j���wJP&S_��������!��@#��|��}~ö8��DيE�k�c����
8͆�6+�߳� S��]��Y4���!��<{�OO�jʰ����w�C��R{�l�h���e�V �|+@�B�ʐ Ur��9b/ﾜCj�-\،��, 8H�zv�Le�_����hE�H≓O��(f�H�@p�RO��q�To���C������������4�#?wW�6�������(-��\N+��C�81�e������f��b��P��us��kQ���|0�C�!;�X֚�["���{C��P�>3,�����IS ���6Ŏp��]	ۄ���o S0qR�MF1͔.��]����s�U�c�+�i������J) ���NM5:d����;]�{<�*S�n��i�	�vfC4M��a���R ~�/����
��I]@`�O\f
�5�\�<��,}���P�[�nq�2i!�Q��9)���0�/R�Y0VV����R�Q@C�v��&�e
��}�8*��*1{3=�a�1hRw�Q�:h���WT�@�5�⮭SM��@�
�C]��3����Itt��Yma�M��Mo�>{���D�q+��rޚn�7�-G���n�P�[VX�5��>y�h��>A��E�11pY��fOv��_aM�T�s�A�T"��������~����Y+�q>T䝈}���_������9�u�*㪹3�,�9�k"��:�\h�d�Z5��F�vZ�Ċco����͏�Ug'~�����h��a��#�E�~*5*Jk[�����Od�+���o�C鹷�RK��F����D�ݰ4|EaQ:��N��*��r漿��Εg�"u-�tU�V=i,cE=�%"��������;H�=��6�zI�P��?�&���5��	�U[��q8w[-�m�a1�5MVeq.�7�	�����<�D1��<Un�A)U��/�1o0|��ۼǥ}�k!���&��-�S�Z�Mܝ&1'������#�~QE��Md�FoW|K]��P��VQ����V�দhq����`��1�x����eU�.�"�2�r)����DΒ����j�@��ۡn`��k�/R���B^(�>�5.[��a��%��-�!|e�1�ʺ�c����e�iR��V+����[��_tb��?�9Q�?�,��N�1�Q2W��`��XP�U��y���Q\�S��lˣ�0�[��ȟ(��FD��<I���딣{�?��WȂ��v�N��ʫ�Z�cK�G �����2ܥ-�t��h�~�_ɦaa���]�[��g����L��ɲ恗%MB�p�KQ.��=*x��y{'��Z��j�C�M�Q�B�ʸOF�[���6�D�u�|��G-���Y�{a�"�x��37j�y8&�#h��Y��{W��S'��b��x=K�F* �KT����s�ƈI��8L��ZR[�Ѩ���h����5�	�
N�A���7������G��t켱��Ǩ�hJ����-�&�r;���-۩{%ʋ�$�f-�"Λoq9N�iqz�c{�k(�i�<L	����9��»���H^�mr��[�O���o���W9����B ���}(���h��u+���+�WJ�P@+�hf��9t��ł����{�������׵V�2��鮶9Ä^P�#Sh��(�XZ�o��ww?ø�Dp;MZŬ��"��7v�"�i�O|�,4��y�'Z��`��3%���"���p��Y��p\m��H�[f�mfm�I�Q+�z�PTzb5�^�/���G��͏�b�X��7�J�sj�顊�f�z!蒼�\Ŷ"�v��9��뽍�p!�{������J�v�j
�[����O��s�N���Co_����y�!�(��Y�要
1����ZZ݅�ɉ�y�GBJ.�z��b��n#�hӽ߂%�`�q�l6�JZ�� �n�����]�` g�p7�<W[Pޜ��۾�צP�,n;G|��E�7t�:����)%���:5<� �;aZ�y�,�,��u��2�P�E��ߊ͕7���⌌9@���n0ė�ư�8l�s�l�����\$�nv"��*L�N�sҜ�g��#rğ�]���7ڡR
��b�m�;��U�f?�_7��}�|��+}ݛ�-(��������X(߯
nM$Ԋ@������#Y �������J���1�
}��p������n#�]��骶�$�l����]_5q�A�x���;/���� QQ�H$������}�ݟ.�#����%��	B�%1%�D>�PS˛I&��腡I�R��t:�mh�KN>���_0���vKS>N��r�� ���K����X|�p��z��a�l�ɭ|��`�(܅�M��i3|i��}5�>Lz��J��<��-���V�|9V��zB��hջ�7fSe�\V����{�ֽR���h���רZ>Mj���b���=�kS<^O>/�c�d�b�%���לI��Jb��sSZL�.\��7�_�A�����H��G(�ƴ>"(Z̿���I9�3C(6�Qbƻ����L�+���"�	�R�e�.���#�sPBFb�զ6�����QqMS������uQ��M���;���'_�x^�������cK�'���?�J>)rc�Ǵ*(d����53����F�J�GNM�;5cA��;~,�H8��~ط��-�_��M�Ml��d�
ﱵ{�<�=�]EG�&.������r���I���F�+�J��R�����z�W���$����E�&�7�낪�]����ೠF���F#�~c�E�����5d"U�$��z ��t��_��YѱΛڲ�
%�}=�
�4�9��24�B��Ĺw�v���%��XO�<��9�K�)����[�z@��_�����΍� !���Jz�}�aN6�u=����N"�hz�J\�EO�J�W'Qy�5jC/Ē"T�LeM%'���y^���1e�G�mD���g�"rk"�+��N�.@d���t��+.T�鋳~0Tak�GNx�y��O�S�]��?	^��A��:��{��� �-VG�p.�/��b���>+g�%������Q�Ӯ�ty���՝
U�&;��/5!�հ0P|o���`�!>�UB�-/�y�.k��@Pm3����H�}�uM1.�KЯ�SԷ����E�Dz2��m����� n9��0%� �)f�)9�#��������W���}�G��[3j��l��$��ˢ�&ش����uez$��(�ɤ�f�'�����G�猙��kG�O#�p<k��B"��q�l�YB�K�1<cxHg3?9��-}�A(4Ǚ�Y�߮��0���[����X,z�SM�;i)�� (!��T{��ʗ��=X©�	��/9t�*.$��Ye�M�O�y��P.��U���^�(\8������� ��16�*v��)�Y���&M.^=���װ��o��r�(��E��`�{��=d���G�&f
ּ�Yh3�x�)��=@�ւ�jcI�Uy4�� |
����9� G[������ ����XlxVHYEB    fa00    1e20k�o�xF���},�Y���Ѓh��=!f0]7�����)|����J��ȣ�l?���N�?�$�~�&5Oz�g ��f`�]?�yߨ�y�^3'���B(���^(A������؀_lZ(�R��H�z��[~&��Jֿl_e�L�p�~ߞ�YKY���6%���9|B앿9�w`jB8oٸ���� 
��71B��D����n��f��
r)����%����,�*��Z�F���X^�X���+�./���T�~��eg�� ]�qD��~b`��D��������ľ�z嬒�6�@B��YN��k��bM�]8��I�흌�h����������嵅�;l3B�o�-�ݒ�X0�@
w��M�Wʙ�\�q��X���g����\�?٤<��?g�V����׉5OU����Gd�~B�����xհ�*�T]5�#�&!Jj6�Ga�������{�F�Qy�o�>��2]:��:ܑ�v'��	SV�U���?O����ĺ�P�Ԏ0��W%Om��� 6S��<�DP�dk٭m��~w��Qь�ǽu�	�'�4D��٬_��m���ɦ���V&'��U�7��3f��:ux>���	�ສk/!�b�Iݔ�=��	�����)e�x�NN���p�4�<W\l� �B �㜵�t���2�M�����xZy�[[1�Iw�ϙ,�VE+�s�Bl�¯�����o��� �d�6M�]�S]b!o�{���;�b07�Ģ+K�r�r�������یC$�c�� Mx����	�/Ϝ�XO�a'�7W��FF|MK���)v~,��K���d\!;�sEKBE�)�4�Ac�EՊ��T/9�H��v�ST1IW@��t�i�E����g.טO�`�bk���&�3���3w�j3�����k�脴Bmx��q�i@�*�*�0+GG��m˱E\��xfNծ����!M�/��6*���;����`�"���tƏ�ږ�M˳�+ FK����B�_빞d���.]5/Fԅ�}'��C�{# �.�F�dq��`0���5�Y��u�p�0E�=�N�zD�`.h��%?��� c�rf��w�s9�q,��_+6��@�dH��+CS�:R�k(��p|/��-x˻�Eb���/�7p��Q�H `V�ԏ��y�mP�<V���=&U`l�1t���e��Б'7|���B�6$>�i�%�ejh��uؙQթj�5"�伇������{� 9/�������W�f#w�Հ�{�l��h�����ܦP;�
�w��O�{i�b'�O2-�[J �yz˽�qY��jF*�́\�VؔC�5��TN}�zyl����A|����T����z�����0��0�VT[E����A�c�kP����`+K~]�ad���U��J�2�����JPy��V;A5����D��We�0��"T��H���T�~���QR�n�ﳧ����GH�A|�B�g�p[�&��0Xm"�+V{�Σ�䔜���j|d�v��ǈW=ڕ֓����é��?<�n[�7*q��ﾴP�ƛ�1����p���;�͍ͦ��y��*��-7 �7��ǧ	���`̡ॉ#�eAN?�|W�m���e��ˢc���jdL�8��i��I����(HUF�*�x��[ȪЄ� �U���N-�п�	Zn�i�U��X˔e<��j��9)�<�;gڡ�#�)�t���O�M�{�@�.P�2]'��ŢZ�6mATgŷ4��iX�/*P-�wf��*���7Ti��
4_@`у�(��Pw�*'`ø�����Gڟ�s�vP�y����5�E��ڂ��k�'�
t���!��jB��n݈�y�=�9�'F���~�6����,��� �)_���&#I:��&X����A�����w�p���nK��r�����g��_�Q$P�ѝ�Dbls#yd5`68�-rg����<��<��Z(���t�F-�8�Z#���Ǟ����ʧ�SC��DӘğ�a'gTA�`�+���xM;5E(��0�$j����z,��a�@��"\�+�p��=�c�"�4P��^A(��+�I�}�w�!��p����3��[[��R���l��&F	a����NCRz��1~��1�w0+�@�ܪ����<��5�Q��:p��I�S\
ِ�b3/�gP�I!�Ra
f��+�H�~a,X��#!�bJTP�(Nv�eZ�-/��v�!Zj;8z*�o[�A,���Sp�зm���F�:�/����X���7��=o�*\�o�ͅ��T�t�G���D`f�m��,w�Ӄ��`iV��oWU����	�izx�f3>Q
_P2�ۊ	� �����?�诲��l WۗÇ�������/C��^u{��<�z���&.%�����|V��^����W��0[�/���*'�:0����(�F����vΡ���������'�J���.H�����ຬ�F�ڽ6Y!&u	W��?3(X��f�h�B���l_, ]kh����Fpi7�Ud����R}���=ZR��O*�Z�y�;�/V��t�)/���?6
��|�}��{���$.����R����&�8�Sk���i�8�)���#�d�R2������w�i�·�(�02��vLX�x��FZQ�(���U������C�1�$�Yyb�@�E4�ͱ>V�{!wo��t���I ���H����k�d� =+N�e�2�S���uo�����VD�J���048�A!���	~�
w�V
g��x�TMH�����ߧ":��[��ߐ�^\���H��f��E�e��S�;���G�QC��W�P_H���셤�	�n��V��}?M�!�����k聊 �ݼH7ѽ�\%Ӥ�4"��e�n��� �x)�13��Q��R$0��ce����0����x�Qt��Z/[r��\d�t�͞�Y�SFF��I=�	����a�h��ܗ,���q?$kM��Y�p0���%_��3R�3�5��eFz[�;:��a���{Go��ҰL���;��ݱk��%U�{�����#M��[l�{�t�>틫[
M�$���WS�iL��hk��Y͓LY?srIN�L��+�T�2rKǙ�a頉ʁ�h�F�F8Th*q�n�[�h}A#`���ra����\Z6�k�ӵ	�K�^M@W)W�"�]D\������

b�"��k�������&pB�u1��YSjgd�o4�1f�&;�[ �N|�(��h�j�X�����B�4$n�Dq���M�����7�g"��mql���ҔBL].�BB,�xW�<g?u��d�+�Y(�/���Ռ	����a|��fg�D�K����%DN77A��N$w]�Y��VL�	ʲE��#������P��)9��Ȁ�T>�,J뇦o����nc���產��c#cdB&���_���Q��L���x��G$��}VՏW[NZ���Z��"�_)ʏ��R�8$�J!Ӄ��9�Pu��j�!�������P/��d�ew!�����������T���J��@5�8�Gw��M���M���q�hV\��!�V��@�q/����ZJ���Q�i1y�GӀt_>�Y̿���C�^���jSf���Gǲ�V�v{(��æ
3w�u �D��� `.1j<��@��c�O��/��fCr����Pq4�!3���yq,p[�xjXI��&&��� n�S�T
��N{Z�9�c�Z^t����D&�rp 7\F�e��g�����t�J�����b��:�����=!5���MK��3ɵ
�d}�nZ���x	D������H�ޘߜ��e�#�r��C;G7zs���ܛCM�veuH��/�uz� ou��-���G��/ݜq�_��g9nq1�4��n~��Ǉ�DW� ���ʔ!.����3�5���t�2}��v�V�]Bmҍ�FC,Q�"�_���L��V~؆=��>=ڲ����5��-afB�$��iO��t�FP o�Ԃ9G3�a��`�D��9�\w��2���Q;�_GbaO3���U��$ӯ��:kȶ�d;'`
S�1�=9�Z[�(!Ĳy��|��~���}H����Lb��մ4��gj�x�L�u��/�+A"l`#�h@2�J�M�����o*�2!o�1�XYG��q����v�hb����Wh���(O�rE��̗�p�!m`��B�+��Q��>���ן�ص���?�`X �/��PJ)N0U�je4�ò��Ϯo�0q���!*�m�o�Jp���t�����f[� ˼S�w� ,(�{����}/&�U�����B�J�Us"�q}Q?Ja뒐4r-�!�+v:��T�3 ��w�i^�����������AvF֓rWa��z:<�d}��2�{堈"?;s�����
v500�`�1��2�ё�ŎJ��n'��jYU��k��i7I��k��n3E��x���,th��N;�7�����Kg�*���VUU���z	+ȁ>mB# �Q�.�K�?�Q��e�ݔ��%Z�!�|O����h l.����w�֨}�.�Z<M���S�wpF��l�D'Md1���!��,�D4M�5N�=(�~ǘb�v."�b%�ǉ�Q�K���#N����Dg#�LU���6bOi�8��������/k��ߜ�!.����xg�8	�$���6���H6��^��|�)��ߴL�=���'Mr'��X\(�*T��1c����J`df�8HR�m~EM>(�XPiѸ/�'שK䷜=�.�B���_�޼ޠH&�s��7�7Sy��T�3&	�����|/`� `W�>�Ya�I	���i�����CqH��
=]$�b��w[u,�M~��w���1rx�������i��d�����F��
f2 \a�0�VHESX���808S������FOy7�l�����K�E+�P
�[/�˂�rݙ� Ǿdi���t=���p0?[��Lu����V��"���,Ҋ 9�.����K^�0	��4P� �ަ:�lLm�~7Y7��h���H�x�z��n�2l��<e���40�����pe7J��b'02���c��Q@��=�*E<�iCs�Cae#��s�IF.<�-���b�c%�x&�r�ְ⮇D��v{6����X7�G��i�B�R��N�w8��Gk>Vw,�mD�w/���#��p����U��D[i�u|�u�\;��!�Hc^�4j@:�	_�����GW�&������ᚰ
M�@kc����(������HU.o,�m�E��GP�vY��ϒ��ixӪl9���A��3�O��{�Wz�Zԫ�5��7�'�%�����"2�zu_fNKۨ��.*���=�b��ʞ��N߫>�20��(�4�Uܣ�;C�$�L4>���Lc*��?�n[��V����1���� ����\RO3�e[�05�Sˠ�my#<E%@۟�}d����(�J�;[���Tv���/��q:�N<�Fi��F,�M��Y(Mx2��C�B��e6���Pi�}ϠB'�����A���=1f���T��b�w&��-^Y�4�c �T�`}B%jMZ��=Pgi�kTQ�����*�ų��~��u$
�+���LJ��0^m/�%�@\ +�����|�@�;Lс P���b�q���EH�-8[	<W�{��w*d������^�s���R�h��?�*�;��6.�=����ތn�����g���d2�������p	�W"�ӥG߮yqN���C���%��FѝUH�<O�e����v-��N�$�u�o�=������k�r���ο�]��%�?�@�/���EL0��1���-}��pi,��:��<�Z��bA��_9��,B�ǰq�P#|�+
�<��!���{������y{=�$Q���tʬ�������;��
x;����������ׄ�b3��> ��!O��#	L�M�r>������݌��Գ�;����ķ\t��y�d��Ql�Gǘ5k�����Z�Nťl�8��+?{�"C�����������n�ruǼ�����~<�}�{I��<:���qSh����Rmh��@�VX�nI�(�^|��n�Ƶ_��p�f�Z�e�Ga�8��@�����8��V�vx�m�y<ǭo!|��u���9:�6fm�տ� ?�f1)�������0W�����;�w�wcY�!3p��4$���D��J��u�ؼ���0��x��q��-�oE�n���eU�� nI���J��0o����(�s�[X�v�
�e��2�$��������LT����7GNy�-��֏n1��<}�e)��d�b�Ϧ�1�U�m�^�M�;tʛF�3�1���i���H��W7J^�~���Yg��.
F�ۦK瞹B�����D��������kq �괈�+>���i�(D�} �
A�{-����#�U"���Ǌ��!I��^�\���47��}vM_��1)|�����Ơ��s��j�ʋJv�d���'���~a�O�?��N�� 1 \�-J��U1/@�}�"!��*�2���q6�-A*Y `�e�Ё�$�,p鹫�`ւ�mA�,gKEzs807ӚNf*�*:��/@Zq;�a}4`����&0�:0�R��{E,k�Ri�� ��tA�����S��!�?tM敺XC 6����I��hŲ��i� ���M�"^/�rl�ࢸ~a��pB�z�g0�G�
�g�-�-o����o*-�)�$��V��0�E��c�h�Z�X�����ɓ�?*EG�F��.�	�N.Y��M���������?� 	�A-E�p�"9ͣ��1���&�\/�4I��p���'�1� ��-����U5jn��;��<[�/�s�U����q�`<�z�d]u_��&+�~�'��E[�lg?�U������4E5AEV:E�H��Ÿ�h"��?̛���8*u�cj����Uۆ`2�	-Ī�`D�MLgY�������xEM�ee�x�\B-�{���cY�b��OF�_\�nh������wڬ��8Ơ�meV>���o�w�����9>�y��u��T�����˚���<1xBlw��p�Y��P�h�5y
Y����:IA�G�Z���%4��7<�v }@��Z��U� 5�y` (6��lw��JM��j�[�^�M?��ce��:G!��1_}B8�|�p�bz��?��v�<!�P����d*�W�
�n_(౶�����k�r��xͥ����Y�<(�.T�y�MRӽ��W����xz=����8���g�gs��5������xRc���39^>�}��)W��5yќ\�}4}�˫�ޙ��̀�X�{+�"�l,ע}��U�f�>�ȣ�[�����_!�i�;�[Y΂3&��
�欁3?��c��tA/���zl>*`5o�!��Ł�xW�i�8=,�?cՏ6vc��[��|`����);T0b<þc��I7j�܄�4��)��K��%��ކ����D����Ij/�65�bc�"j*���57�\uҝ	�	�����)�y�>AE8�f4:	{�Y�D����XlxVHYEB    fa00    1e50�5�J��aq=���W�O[F�p����r���������]<L#�Y�>�0Kƾڮ��d	�Dj�M�@2$�1�'�k�>b)(s�d�j�V��n'<���)@tH������� �³�%���)դ:�'���e�IF�&[t��O`�jf��Ǯse�8����M�񙟩2�ȯ�"��a�K'jy���OM;��ːR��x�����E칕�3���� �!СYzA�aqC�w7�Y��IQ�����4g��J$V��p�41pN����=!bY��-R��&��!��r�pCҧy������Մ-�K��[���#�T%B����[�/�cAFH#��qPԐ[�v�g�YP�O��BL+�F���3R[���8��5Iu�!6#/���iL���C�@��Ϫ���/fܩ�P|v�w.��<���F�ZN���xx%����]�����.�r�}��/"�F�X7��f�p�MA*	�ďz��f��
\"�i_܎
8p�ξ�H)�>�sfȾwX��%	J2î�����½PJ��P;]��3F@��P�7���g�Y�l����������^&�* �yU��W����݅�ܢL0�֞*L����Nw�����>λq�������,���]�����6 ��`�?z�Y&.�=r>�l`7��_V�"�f���)6�+���� _��T��-m�h�ljy�Jޣ��>�xx�k���'����	�+��Υ����0��X��T��eRԫ5TQ�SQ�H�Z�*���r��>���X��=�S��� �EY�T�ro�B�d��R�&�F��Ϧ�ti�#��<Bf��g����9�)~��6�7z�Ԓgذ�'�f��R2Ta,���(�/�2A<d_��x�,A�����,\~���rozk����1T�&h�q@��%��1��ŴmN��f����J����ܜ%B��ӆHS�ת&km��"�8�z�8���-�c��=��N�^GH� l�8?�h�^D͔��A�]�겏������f���'����0�UP��'�qgGZϝ2��B�!�{�ө�WS���.=UV��(+���]�B�LH'X"�����	��hA�ACTx\B� ��>�ޅ���.F�i���i��S�����ٶ"A��vb(����8�5�� D�q˥d���t��_y�����)E+V��Õ4���j�i�"�����!����Ά�2�Sø���DB[~���>�#�y�<��䊫`2�~%*��Q�[u�SD���KƤ��k��LQ�UQG!��5���)����e6}�U�w��|�Y�@��Ѿhv.���Y�"�D�@e��s;C�79��E���}��!�E�=㸅[�����x��Z����X�����T�_ �\K��ꯈcHwӶݽʷ;�Q�y����V�����ɹp����b�ECה��.Ɂ:�P �F�"8
�C�`��n3p��|��ޚ�	Zo�����=`��u�'��]��

k坈S�2�,��բ���Ȣ���e3?F��:Ԣ�x�F@V>&�[�%<���Q��+���u���v���miF��n�I
�V�9�剬CPМe9*� ըa�H�G��V�ͼ,$��9�T�B��)��[gj� �ce���al�&	��z����\ΖL�ֲ�jƠR�*[�}�J��0 �͔e-��YO��QC���b�o�}&�2~Ά�9e�l�-A��H������/O�CWs�26�1��Ϡgi��Bۋ��ڂY�{���<�Ll�mT=�+��|��u|z�~x4cQ�S`��Ҏ������N`U�ֻ+n*s�R�������-�o�5y�̂dH�kL�=+��ŲY�B�Oq���1�eS���y��&x�D���U:}���`�[˜�.��Tr���^c�t���lT�p5�{�o �N��3�1�+�0�6�h7�Z_n��{��7��؈4s$�.�B�M��9 �(?C��i�0�[;H�M��{3'��ak�()u�1�v~R�/<�0�|���#�]<aq;������n6��'�����	9��z��(G���N�*�rG�#Wc?N�ſ� �>C
��X_;��~���c�V�a�q�?3E@(���(�T��緹ā=�D�@�2��3.I��i��1�j��
�Ŏ�O����e��h�&[E��yEךT������~�#~*�gjŁ�p拏"��E�z&�u�;t�h�����5�>�
ۣ��{��[���4�ʲ��4�F#x֯��z��
����<�m\��:KH��nlK��W6ԯ��k�f�!���fi�ʍ��1��V��N�l�.����X�'�����wk��^΃W�J�_�9������2C�s�ߜ�����>EE]��+v��0�j�IE�'�$����Z�
>�,\��6:��#$ޅ�:��A\���
%.��d{P9jH(O�=�a�֏CM����� �5ڲp��w��Ɓ�F/z�*��sE՚��:,M�i��c��}��L���:^�?r�P1=���D��Q}���iG�=C5R��}7�����h�J���;�`���m&L�Z�5[z򉪤h�t����$�ӎ>-hk���R(�[�;��^� ��k��@�����Bq!��ևU/��4�Tnp�>����ȵ�����)q��Ԉ������1ӠP9p�Om�1��N�4� ����	<@+�Z��{����>][�W����k��'��% /����(3vY���G�� �R	똏�K�?q7�]��m �]�!��7�Ȟ�E-6��A`��
�:�'�]ce��;J�tJ���C��uB��]{\zG�?j�;��9��� @� a���ʼӄ���a���w`Rʢ?՘Ai� |W����\��L�?�Rwp��P�p'��v�j���Ux�����<v	��/{}�~;ȸUIj�J �6�D��:�ݜ<EI��!��#QA�xe�Z��k泹ҫE"��lE#�>\9�.dN|�s�ɡkT����[��^֧��8C���#��+Oij����}�T��0]�S��e�*��W�FY�Q��� ��&Z�*�5�S7PI�o�'�ۜ���ı�����\�{|����g���՟��v��B�$�=���;g����վO�v�~|
�����Q��u����}����Ц�"�yz�p�6����?��W��=.G�ȵ~���ueؑԇ�@�ߛ����ŢrF!kMh���2%�IR�o?�8�o�b�=ٜ�̶�G���:.8�-MM>ѪA��RF� l(h��S�ˬ��%�Es�36����T�&�Yys��|4���0Z�z���C\���TB+e��*`<��.���L�.s�es�BL{��k�T�������?_*��l�HCo↱?����4�`=�E9�]��}4�y+|�i.
��%9�@S8C�vf�ʯ�o��֪.ޘ N��:?�-Jԛ,]Ut,w`p��� ��}�u=��p,Z�s�r���~;�e���K2�zo��R㤕+is�h,@���7���	';�On��\F}Rn_�r9��>��Zz��۶��tB�M����`�Q�'�<�`�,E�Z�;�7~��B,��:��V�?>ܔ���������g<� er��)���8~�YPk��C�V� S�2�%��'�\p��t��/R���o�o��0��Xg��;a�
j��z�E�c��R�*��ġݠ)Qt�ߟ@n��5���:��K��g�?��e���ݥ	�,�Ŧ
�S���;�1��"'�]/����R����|5+d�I�ؤ���t���_()�t�������Y���)f��ϒ�\�B#(���s�H��,�>��<׿΁:S|i?9�ґԶ�`�y²6<׍�c�d,0�I�xw5(0r�fǒ�^����?�>ũv�f�'H��Mi�rʋ$8v�c��R:�P������@$�`tΉ�Xi�c8Q�,��s��+�|'�z��g��K0o����Y�`r���$s�Fە�\�>,ݧ`�H��~������͕�����Ay��h��r�ޓ��w�턷�.<�p��c�4St��17	�E�$Z&j�y��!��7`���m���%	�e�脙鵬���b>$�TM��l���I}�Z�ȸ:Y`�o �|��� ������D�����j3��Q�1/�Hj9\;�F��t���z9�jt`�oP��4���Du�p�'U�P�P.V�;�l��5����'Z��KL��:ѷo�k��֊E�>^L�kI��] տ7ǘ3�)�_��Vz��	��]��2�I%���Z�Q�@�U�I"���fə���k�`��!�,�]�.Eh����/,�nQa�a��d�S��Fzo��W9�����7J<���Y`�<�ޱ��*_�6�������jr�Z�D���;J�Q�}瀰�a���ܿ�l|f�����)�|����e�G3�l��p6d0c�Y�`��L՜���Jc?2�&�ӤBA��4>�r��_t �i��Ì�0tzD\H��,[�	��&f�X��R �Z��_ӼJ B���0���.�R8��NL�W_ń2J�������%ì���{�3'vC����n�^�Z<�6H�J
�.�P���BC������5w�
��T�Y�0�=AJ�4a�F�R  ڂ�(H�ǏQ��/3���\��g�
`ҧEe�����1��%��y�z���;::�2�6r�؁fac�鞔��Q��T�Y|t���1
H�,��8��z�6w�
z�5Q�W�O�� ��⣮!�GA}�����[[�a�����!��׶���Yr�-U����Ҹ2�������|�VR%�]��7��W�/V��\A���%������������LA�͘�TW����U(���B��d�mP������,f6��m����Kbᮇ`�΁��G0��
=�e�J�H#��/ ���R��?*�v�M�Zo�c;��E�?�D�1�EyE�,6��M#t�UNT-�A��[9����5�T1���W<SFB��>�<�!�GGl2'Q��>;���V
U��#�|�ha�����oM�|y�*��[/\�dp������ϯ��vȿ�m4�d�q����\�z7բ��%�#OWT�.bSt���0-����_TH1���4vl��9\Yo�vUC���lԪ-�x������d�U�ckﺌ}!�Xò���3,��5�Qi��O�����g�����q!�n��v. ���OJ��m�4y�[�L��C�QC�F�rπ����W ��~�䱈��h���l�=&�S}M��<�A˴�o"�;��C�ۮ�j
�돘.*�S�1������5Z$Z��ʢ~ϓ}�F����3j�ӌ�:�Z�neR�%.4I��G>(1zv���!ԅ^{��˾����>�i�(�="���ۑ�,h�b�v�`:�Pg>k���(����y��R��1�"�O�u����$Q����00��|��&��$3��"�n��s�����t�G\)])��v�-v'@M��Z������t�I˪�3��x?~JRIm}�������Vס��ޫ1��CN��Âd� =hCE[�0ND� �9���kW5K�X�,<_���0ۭ^]�� �Wi. l��%%����3Y�ߓ���_CB�6�_� Gx���H�6��(����O�ؚ8�Df���v�	���ϥ���Z z��F��%���@��?"�㓹`����c^��)��j��йw�&�iJ�#�Ԉ��t5�6��#͇M��K"���3B[r9�예�<%Y���������1Tf4�C�&��U'쪰����Xӻ�T�񀃨߻���,}u3h���m�:�P�_<���� �:���[��i甛�vBq'�*��(����L_�u��?m�ָT�K����-����4��6�%���AHn���;��S����]�U��Y��8��H�LM�[�B�}6nn��[@l�ѷ�ń�N�j3v�O[ƍ'�e�_2��B�{_�D@�/�#:|?����&��f��< 襂�y�8nm1)��!����%s^n�`"�\EI��#/���t"̤�+�t���J�~r�,0�ӁS��	^g6Et��FV
�t
���Z#�5�a�t���������xJ�C��8[�q�JG%b�_\���{���뚶���U�O(�{��]S󫳧*�ݛT-��9c��!sx����+(l(�Zp�v�ѫ='_����T���c4�d��.��MB�C!�ܭ��;ݨش̭�V[L�.=VU��o��� s0�
�>�P�{|-
� pd�6��":���|e�L$7�3@�E3c��\�D�!R��:��T�hg=OiJg߭����KIhͭА�m���󉞲��r�_���=���A��vb�?<S{����xP���Z�&�&�y>��5��"=l�
��\*��)fu���v���Yߤ�¢���ܕ(�6Β�Ĉ��{�M�Dݝ��\��:y�������D9�~L+?]�Kn缒�Wڋ�J�^���꣯q+p��9��	n4M�lT�o=� �=�[X#	�����ú�D����p��	�B���"�t�{�=h�����,�M&��zή5�?��(���p��,9��a��`���l�j��";��K��u����t����t7ߣ���D��&*�2��wr�؛��e��O�8��֮hz�9\�Rr�3�5;�wf�� QV�G@��A�J)Y)f0�+�^�:�-�����!�f��|�U��Л������N��[v<	�&���ۖ�1��g�VlW��j�{�Y4�@�2) �����u b)N{i�:΍3;Ǜ'��~��x�tx�@(�P#h��'��5�筋��G��
k-P�����D3%����^�M(�'O-)�x(�h�p��QZ ���C��e_���d�[|ͦ����۬c��yJ9�ߙ�x �O��)!@SI~DY Hd�Ҝ��^eX�k�0͒̒+%�|�|����N���0�AM���{�h�\8]�h�Y+�����l_���48/�15H�Q0�R��<� }�g{{�Q~���� ��<���h*�2��rv!�a�k��eVX�5�m�v�q[n�:Q"i������ql�j�
�e���gr�'	X���W�#�9�k)ʃ%-��pi�G�_�"��7E? ��^sU����ӻ_-E1��/���U�	����X��:I;������rQ��A�+��',�M�f����v�$�p�\���+�3�3��§���T+��Cw&N%�Չ��x&\��8i���l+�0M�#ԁFuZ�X���Q�À�'��c���WGNQ���M���+cӈEe9�U,8=�ܸ�,n��	m��B��?��6�F����b܊W�&S����X�	"X�'k�3�y^���S��d(d�4�36���Wʾ��51p��@ �*k�X�/���� ��s�h�u�(\0N[�G���bFx,��s��HѢ6bk�N����[��p�}������G�֚�&�E�E��q�})c�OVp=>@��:__o�.��H���Hm8��p��5Z.���3��?lXlxVHYEB    fa00    1da0CK>�%�ٱ��`s�2�د)��0�3:��=�Y�Y*+�i�����;�cP��~� ���v���k3��\�������Y��/Qw�s�"e�R�K���*T`�D��7F��n@��+w�������u�W�q��1ql;l����;��~M�l��$q
A�*�VNu�,(�o9aRj��]R4ik���J5 �x��uЎ�P������l���]����������@����J0d�o'f��o�i�1�i��CƲ�侯+�Y/~�b�Ϥ}г���E}w߈�ʯw Ts�Ǳ#y{f��g'�W� �	d�M�G\�O�:�`P�q�缯�]����<��1�ԥ�o�2�VJ�(�ñ���@jgu�/\�̮Ce�Z�5�BB�	��!	�c�z�7�����9	��(_`��bfV��^�~���t{���R�Qd�/�v�@Y1L���Z yP,�cS�O�t�CZ�sT)��� 3��ύ>@d��~��'��oVI��@�(N�'D�[Ԣ�4��Py"ވ�~��	i��8DZE�����.��L�N8��	<�?�;@w��w�x�O.�k�6w���u�Pi�<B;��K;a��j����83Z�;�{4����ޯ���9cJ�c�ߓ�� �-kMJ��I�rO�5=��:����{��eF��.+5^Ct�قDAHH�ؘu7_t�d���?�M�q� �{]e
[?q��D;�x�,>�fP7��K�V�`=7ρk��Mۋ����o���K�7��DV�rם]H�w'��/�2�����6����U��'�Bos� �9@�/���)�:��J*�4��F�O��c�/6�/J��������o!ȋm�c�tZV�I�dJ�jo��\z��c���R\F��F��$Qo�ٌ!dZ�b.T`��z6oV3������@#Y�l;�"]q!�Zv��H�L��"	ʖ�:"�	�C�!�v��x�����t-3`�T[nt��PA�v�޾M����������MX���i넿tٱ�c4�׵��3!�(���`!�eZ�F��<jޒ!�'س��lYm��@=*�lHl2j#�PlD</)t^��p�$��0DRYT�ه�D����������M�+�����j�&�
�1�+�<��7����*��E��#\���%#R�<�1)�t����|�ἦ�Ag�]�:a�
�S?_�S�~��_��i�ǝ�eߩz ��֕��"y������Ԍb	��|�3`�8~/���v�(ܺ� c����;PB��~.��E����*��!a��0����%ʌ�@��Z	r�98���Jn�&�+-���̠�ۃ�L��]����`PY+)�R�7��I�q��I,��ҧ-�T�r�p�b`�̕X���)5?��S������3�S����c���Y�z����ߒ�ϻ��D&ঀ����~�k�v�G)T��qF�F"� 3뙰ڑ\�n���w�#��[�g|��'��:c�k9�̗c�������L��.9���b�g�6R�hT��²W�s�M�J��"���)�]t���B���f����J������h���QM�6�}�=��u�txh���j����y|����dVV�'=hT�1��1��g��8d�;j����Ű<Ɣ�-�E9Å{�wEop�� �h#N��1�V)�\�\�km_��[D�ا�;=�ڏ�l뵖���9k4̩b�g?͞�*q���@K>|P�S�p��̑bk)�W�?@-�F���&(�#x/Ɵ���.������]���������%R��zДU���"�+�!����ȧ���!����>
�,a๳ק�@��2����
�<���ڄ�3s��gWdt2���Kx?�0�ښ�g"x]L��������6`v4	����dr���y�	��k㜋���A�U �q�;�Sғ1���0�����޿��y�?�@��Oq� ��7s����G���\y����e��������41F���?�.?��ɲ�\ص���'�? �Η�ú�꼣�SVJWY������օXzF�>Yo*�Cy�'��lAD��?��Lin�)�)f�����2R�;�!*VI�Y�7j;x����.���F��.��v��!sj�.�Vң�1MA%�NSp�F��p�ȳ���ۣ����o��r �P�|$��*�Qn�o��e�'�ag��O�]�9=���������2�T�@S�z�އ+G@-�[��O��7��,�ލP!�#���3��P��Q���S	����v�۝��%���k \	:r�������Z��J^$QrOå��K'~�����(`̧$�	�9�}@h��QY3��kar��%��U�#h᠂��Ù��ڢ��-�$�wԇ0�c������=�)��a��/[p;FoX�HV�S	��^�@�x&�P�Ïd�&�����~��4�w�/�QM=�]X��4xv�yi�
.1�u�e>���|궲��
ς2v1s����.��%��04�mݢC�Z��m8�
q҉�߂U:H>�g�+�x�h�u�3��bg��e|�).�c��	�#���|�7l�����������/����30�X�	��7"nI�M��S#�֢�½���N~��-�oZ�����1���+�J�^��Ԅj��q�E�(\GE�-7�p �By���'=	�3'P�²UF;9B62Q�%��-a/��� ���T,�I#l�z?���Ch�f�8�[�W7r�K���&������lc%��kejs6�@��Y�Y��7���h �&rd���$+�9f!�3>�[b<�S B�t�7��+oy�oa4D/.~����zE�N�������FlD�*1��d����M��(���� ��^����$ڿ����g���z����0@~{�����,+����ˍ�8�HHb-���q�vl�(y�/�ï+�l1�6���y���6�q|=��+Sj���s�u�7�^r�U���;F���u[����3�Z�"�܁�RZ
z!�� [��"���ڸV�d�y<���Tr#u�SP}��<R/n	��R:���g7�����=@�,�����6U_��mҡ	�:���d4o�0z�|K�Z�}������.3��	y�Û��I5c��,w�0
���r�S	�?~�>��q!��{
N<YlN��"��Ut�=8T&1ؗKQ�Zqe�J�Wj��s.]��#
��_~~z���+�^��5<:�I����ۂѹ�A0O1���jZ¬��-K9.���_�����FW-~��Q	7�����c~o2s�.��Y$���F!�!�/���N�t�\�5� <`��h��8ؘ�-9���T�b�O�a�kZjt�G#��{�� 7�5�h�����UҤ����X�3���"Tj�[/Vj��a�Fົ���յ3���MuT��Y{I��b�,%JV�6Y�1��\��j�_��y����
����qI0|N[�܅��9�jz;���.|2�R4S_m\�^����#��9i4�Lφ�"�E�����q�n/�w2=�Tt���[�K�$Z�)��X]�<�WB^3ϹW�Br�\��CH��nv���C�+^<3��f�^�/v.:��q���.�	�\�/�U�:�8�bWe�2����M���N�MP���� ���&���Y��#˶ы~�W>W�����$��g�%�t�r���.j���F��˚ёi���:0Ժ��,z�J_-k���+�TS$��d&���s�J�����E��cXl��U�l$��8 g�e�r0�ޤ
��A4i&�֖%�-�'�GN��h9�������99��`!`�@x7����S���^�Oy�,:F �^�����f�|k��D��sL�U��V�8��C��I����rR�	���s��Ov��$�T$G�����<6m�N@�>�I�vh�$a�w
|�71b�O	��̂V��R��7�m�&�W@�J�6ڡ ���-D�Iw�o�;vqJ����\���h�v筊�1���!=���������)��ͪ2{�D��ۖ�)���u'���%����S����cČ�	/�xZvr���Q����ܟt�IV�t=�R�����Nr�8wQ���2���Z�a�IT7��26���~��V��KU\���%_?�q�� EǨ�А�$*��!��0s�G^v��_C���C�35x�V��e5�\u���Q[Xu�J8Α��]�i�<��N=mg�*y�L]��-w �C� ��ⴲ�s���F�ʭ2��w���X�)�f�,��"�k+X7���爏3ٙ�]6��I���Oy�<�g/�i�L��6���Bѽ��R��B�;�ߥܫQ��C�f�N��]�Sn�x���H�7�I�uĽG,�Pc�/7��o Դ�|�a�
j�/��^��⁊/ZB�~���c�;ɨv,m#j
�Շg��3�?�͕V�	.r(�Q��ӵ��J�������N�dD}!|�k��4�h��rQ�HL2�:M�ȪcR"�C��:5������W�a� 	ݦw8a���R��^�x=g\e�7��RF��H堾}��] X������fQ�J��K	�t,����A(�9&�N�ظ����4 3�=�`�Q�c+H���a˝d<�S�<�Ey���(�E���Ba��;u�SP@�� '��ɰ�߂S~z�d������߸��q���{�JGaF��_�_�a�
��E�B�+'[��czҕ��}ͪ�z(�e`]��)������$��<*T'ah)�0ND[?� �­G����%�9bVO�)��B����
]m�1ܸ%�ΟI.��
����pJro�<���7sh��@@h8�3��ʳK����'4$�hz�t�Hf+��|��O|�8�>+��k�(������P�%9:��O@E�!��T����-"��G�jX�x�XS|8���w�,�E����<��T�ʯ�L��ح���9���S1'aؼ/
���M�u6(���^����O�Ct��'������&	���`=�%}�U�jڿ:���	����,����9זݪΉ*F�)�̌H?a�^�I0�%�ɷ������J��F�E�E#���h�о���D�x����Iͧ��μ�rK��^�G-㏫v~��6{��X2/9n�ʉ��XB��w6����L�4?�{�����R�)��^�T�T���0���?��Q�#�U?cNT	��e��8^�PC]��o���^y�J��C#+���׌�#f����r��IE݉P��!��J�����oG�44����"�=��q�v�t=s����8$�
������z,�������O�~�zp�JGk�i�!�*��:�Y�l��ӿJ�s�����1n#� ~ޛ��gN�,���=!���LRS-��u98�2R���@��\�v��M�!6�|<C���ff�(8M{R̙9��{�L��%i85,_�g����-(�-y��V�
�{�k��U�8����v���y
�j��6�)H��|�>����\zm�ɱC�5��u�rm��{Y�ux�֦\�:6LJ���T1�l���YM8�$w��o����9Q�;mpi��v��j�!���1���Z�e��n�e�A��E$9$���W����S�϶.��y��њ�ǭwR\���X?K����"�������w'!~bl.�sN/�`Ĳ�C_(��"�"��[�Iv���gv��5�#X�sK٨B�\	h@�YFOc�<'�9�>-��&����R��ͱct�vJ6��/Xb�)�o�)`վR�u�4�䎣�z�~�G�^wsh���A٪Dո)x��9�E'_�<�cXCwX�� %�4�ӸD�p4b�q��W��`XZ�Sg��88��:BRU��.�z�����A��!�?k%�p�g�-_��ĭ{ľ�2�����ձ1�c�b=F�1~��ͼ�M� �ՠ��8��Pը�@��ʡ�w�P>}��ŉ�����x(}��<Z_L^�{�h��4���{Q����l��"�4�������=	 ��t 8G�D�Q��D�$[�.6�;���p�r\[&66���
`�C�<m_~pL��.W��ThRL����9y>F��R�c��U�{�ݟ �iU���3QIP�P���-D�`��V��&���ch�P�M�0�It,ҽ#���2�h=�
* ���Jb�Yq�|,�[7�9k��o������ʢ�������6����?#s�Z	^�j+�}F�Η'���pfs`f<�vV��?J���c֗ҙ�>��p��*X��u�P"�>�����Zrw��&KA�m���43`\	Z[��V�pp�5�����{�\��f¸��+��Fap뮢���.8�a���z��䶔W��9 qsŨl(�%MG�"a��|39�����^��wY���P�x�So��2��ƈ?6٘�Z�S%0���q�of����ͽv���`g-�vD�bD�y�&��"�u��('q��p<}0�#R�}�#�UKRRC6���K5��󪯷��!�i*���@���9G��d�\}�urq4&�����}�$��!2'��}a���!��D�:�:�sQ� H�_���N�U����![���x�
�D'!�,�YVE;f��#�.٫�� �)'�<�j���?�ħ@��S�� �=�A�Z~~D����0�6I@��1�2�v=h�3��T����:K��yh��A'2�����h?qC�w˵��丌�X�������P���S8�|�	\4�%��z�u$Jd2R�"?�Ȏ�7s�Svͷt���w hN�U�ӄ��?��WH������*5n@�]	v���Y����9'�G����&\9gBp���{��N��y�T!��o��g�a�R��#uʋ�yQ|����r�}��ʻ�椦8z�N��	b����c"��զow�*g7�̷�p���`C�6\�2k��e�Ɔ��:��I���$���h�$7�6T�.)lV�c�Ig|�G%�FI�⟣�s��QSR�I^�0��S���ȍLGE%��;/1����5���iq8�=uU�fHX����x ëT������2�b����y����n��M��1��Z���:��"Zx�l=E1jv`M��e�XT`A���O��A�qs���tب���
� �s���Y���@AȞ�:!	?�.�ˏ"��v�:���b���$�u�L��ȉ�����4�����_��>~6���8����,��E���D��S�ȋK*�1��}��ҍ��L���u�o�˪�U����HBD�1/��}��_�)����n�/���;@SA�&��،%C�1�a	#��k�~B1�P�,�7��}����p0"�ג�vY^t���.� tDe��O�XlxVHYEB    f314    1b50�W��U���uɱ��Hs&
���9��)�x!�H�&�y�������*~�K�J�[�s����������?�6n�,�7{�l�%>��+�-Q��{U�KŖ���5b!*��/��P?jc�5]b*�h���?����%1$������&�
rDN���5��l�;6wX��ū�T�}N�-R��HZ��Tr�+0�u���R�.�1fM�F,	��]��nkt4�#�'��m'%x������?�Y{������%�B���I��<�o	�؞L��xK>�t9�����v/���XA�=y��G���8��M}b)����
�}���O `:��"��D�^t�T�����+�'��l�dv�,���-�N^�!����Y����Њ�:�q��m=�o�e���?/U�+�S%o��`S��^_��沛�2���ӕ�W9�C�8h8�^���*m����Q�_P7��B{I�%!>紧��&kU�oD��\�P-�mui�L��e��f�_hb_28�����6���6��N��
�q��['�XRsO�Y�ika�_��Eɑѽ�>k;C=(�d*�o��핀4��#�����F1+���3�[��p}t�Aq$��vl���5�"G)?��tY�ACp�V�6+
�0��c���Y(UC��;�7��n�l�7���u*K'�?[�g�7�#��v��o���W�ݠ��Q���Y</ns��r�{[������$�]ѻ����J�Z�FW��b��(ڪ�egw��i�� }��,��V�����ǪEG�U!G�G��.�"�-I�� ;�D��3Zb���?��Ss�,�����������U$���La:�MuS��k�o��޷l�X�r���U��?v/n�%D�b��)�$���S�Ցd1~�"3#YB	��{�<��M���l�h��3g�$s��Yg��EO�W?�RIBF6U��r��
�u뢴��j'�Ǻ���Im�Z2H�(�&#�A�;�����9��H�$�)Ĳ��4T�$��G�|3n�����8���ԵW��6��z��Q���o�̉$�!�7�4�+��D1͏ߖ�..R)k���	;T�`�gX�$w:��r�؝U��}DK�&ڗO�'��E��NX��J���$����΋9.�Q�n7x��˚$z�~����1V���m�oQk�;��w��c�O���	��8*s@جgB�8ї�����cy��j3G?z2�� d�VOk?$c����zk׵���fXM$�6V/��z�nv޿u��-c{�� ��e���izx><��c��9��կ�j�A��F�>���zx��,?��Q�	��b��$���r}g����pjÂ��g��r�M�g��Lh�d��SӮpZr����`�N$Wx� �U�tl���Gr�֯�3@��N�e�8��u��U`/�<�:y冥Ξ��������Ux!1���������Y��Q9<��FQ�v�'�YǸ�q�.ٶ�o��9l�m��#�7�Y�w|<Zt��߰LN;�� ��m�>��<9�aL��� >��:�b��3��B䟆R���bᐎ:��1G:ZxgX�oxzԯj�8�[pu)>�t�xI��-}���`�@�m�*P�glA׺��i��S�����~�~1�t�#��̻W�H��c5C���m+�5(�+����
��?��U!YY���&��59"MFA\��î�4���m��%���|��ǒ�!^��\���9L�e7�J��Cu�^�H�����Yu��-X��1��#'��kZ[���5��3�����j3��]���蓎�A��hFp��Bf���\S������"�s�2�xȟ����;L|R"T$�+�Q[����$���ݝ�J��ۺ(��ܬg��?�bn���E;S��)����B�b�'m:�\�.�Sw�W���.Vﰪ���'~�{����t��3b���^�}`X� ��=q��p߉�����b�3{��B�Gk���՗LR�l�5q�`��2Y��FW��e�J��=�W=��ZS�p���X�/$��#§$}���J
E�@��`q�'U�tn@x���8�b[ш`�6PU�d���$�����M��#�(���\v9y֎�3��y���gb�	m8"�]Wذ*IîD�NsT1�d!f~!�,}�0��0O�+���C�]wT5G6����mn���y.W��R��p%�5�D��d�{Il�It�J؝�����VM"y�m��NMt�0;d�.���/�E�n��_Yg�Z�a#�9�O� %������>%��<P�o��_~K�3F�n��пu�w��jF�Y+��	��U!v
G��bm�|P!"�=m#�@�ǹ��x�6���'o�9Yi颍�q��m��.^��E;G�V#��%ݣ��~�y��#u�L�"o趏2����noH��w�����+d
�})l�~�B��<Y�|��(RH���j��R\��X����� Z����$oJ�QյI������Jv��=��?v�r?~��҅h���o�X���,�����G��s�
a1�Ra?��=��|ra��euѩU�!)�é��ͱ��%��6���n��	������xR�����@Y�W�R�e����Z"#݉�O����Cw��/VA2}��@:QGd:kOl�m���0?�5R����1,S�E�r��:�84�	����j��eZ�s��������Ғ~���@?�\�1o�=#_���nF���&���T�A��yM�@�JZ���JQ�ďY5��G*4����@����U������w��{�0�/���hv�w���-L�O1�b�C%�}>媼)�7�2�n��PS�[�TV�X�f�` � ��%�v�CyC#�5�O�'P���ۦ���I`�]pL@��>�{oqm�����Ӟ!��5N��	���޼��>� �z��aJ� u%8ɦ� �����Z�	���f(��)���֓���x�l�0���T���
d���b�H}N�l6�_�,�q�p�
��_�{�@BW�a hi�s�y�`/�T'.�V/?��D� ���Y;�A�r+6��N4�p��ߗ����?������R�yu��T$s�V��ЮX��ߙ����M�^y�k�9GD�Ӈ�{���Ug���������/���*�{ c�ˁB����	�8 �D�6��o���aͯ����ߪ�[�U����2���ւ�L��aZbPc��*yoL��ð�SqFi��`yᴾݤ�A'@��fBd<�#���Frߟ���q�>������'+;���M�S�.#	F��&�@�K�O��X!аH�og�2Z�
W�:�w�||�8�,`R;u ���V+�*�������((s9�,�n�p��}N!�T0�%�V�i�O�'h�})��Y�\=J.��zj�/��`����Ԣ!c\x��+:(e�C^���ϒ�$�5y����_ԍ��8���/cVPwa�<z	C�,���*f�Э�M5C�J�	���-�����Ȕ�d]�gþ'�'q�g�-#/W�Oq����߲�Q\=�۹�I�

���b>K1�l��+�\/�tZP'.���	ѧ��)�A�Y��Y���v?��@J���n��{��d�08���u��Cx�}�˝ݗ��r���@_��ٳ-�:���t߃O� .H�տ��h����;a׼?J���Ǿtr-��7m"Mk�81MK�FG�Y\!ĺ򒀿�U��\�fm��+;�@�pa�H���<
��8f�W�3b����k��ro3��M]B�y�A�X����i`p��Rϸ��wi+�`��U��L���X �t%lQ���4�6���C�?�
ߒ��}��ع`�B���8����L�/���ǌ@��$����o��	�;+�o[&s��HH��Ӆ7�]�����(E�b�չR��y�S0>��t���_�ѲB(��2(�:��P!�sNʵH�k����輓�R��pS�����xd���PO�7$ꤿ�p�ɻ.lD97�m���M��[��z�s2�����W�"�Y�����zy��h�vfz�+7��ʱ�Q6q�ڂ��l��y�p�fa�
��F�d�B���ݶ�<�҆�i^#�8@�D�l7��=��VYI�6�xx!��1�!�遠�/He�	��f� ���֞011m-x��C�a�����p��5bw������<|t,�n��2ʯ�"�w�UZ9H^�&�oI��5��~��ص�o�r?��r\s�P�j��w�2<6���"Z�j0Wц;��Y�)�N	>ڈԛ�(�|;u�b���*�*X:�]�59A���%�&��(��U�#	�^:�2�|DPg��֙#�8���CN,��rI:�i������E�/�p�_�e�	�1��c�ry�==��u6�H�[ӷp�p>Uv���E\B�3�1���瓎x}�j4e>�;�<&����icF�=W�@��;�7����,��'��#O���Lt��{���h
Cq'�p���\����B^@�O��F0ҭ`�/���ynV�Z5�e�eһ� ��O��q�$8��"��k1��wTA�&b4�K�r��Po6T������rA�Խ:�p6yI2�賈��ox�~y�LT*�H���GR���"wPL��9�{3�W͓c� $��e<����\�T@l�Lmk!h���@�#U�wn>��>ɪ�ZV�Y|��Ed�s�鹁!7�Bi2%w�q�#X���<������O���ܕl�����2bߺ�`ia�9�")C`ލb͝�>��9~��Y|dIׅ�d�e�I[�)ݻ�qr�.d�m}�e��c)-��pL����J=�#�Ou�(�c�L������hl�	�Z�F�#]5�>�<uHh�N�'��m�3[߰H����E��\4�K�Dyx"��H�fE��p�=D�Z�-SΖX�O�NP�����Ȣ�;��ԗD�X�mC��4�Ɂ���������Sk�q��G�kLW ������z�a��LNYw�����kL=%�E�@3&�ո`�Q��L�O$ի~����8���[�g�r��S���R�&Г6�,�-�ŉ�έp`"!�/��.S�}f;���.Z$r0����\�ψO�G��M��#��ۛ�oLS��[�髷/l��y	'�ב0n�=#��~�)�����[��2=*�L�mI!U�42�<�H7�@l!Kj�Z9X��q)<F9|�mYhi��7�]���76���a��IOmi���e��ɫ�&���}�l|K^�cR8k��?����cl8�B�w!}�|_�4�q�cj���#���j+��$��?��@���Z빀��8W�dbF�J=)�����,�@f��&M�7�2[�s�l:��R��"ߍc��zEfl�55%���O2��})4����YWZXh�����ȋ�������w�?�nuaK7����cp�;��&�\�r}�t"��?E�/Mt����<ÿ���P�̀�ת�5���r��HЙ��F�Ӽ�zU ��������;zzz	�pB��Й�_U{���P�E�fYTZ�F�3�'睷����]o�$+\�[�F�bO5^�8Q�(9�����������X������*�J������a�Ӄ�<����%vB�Kg����ț���`�*�0^GI#�A��e���y#�4e��y�7=]�ܗ���G��Ц�K�����<â�Q5a}^y����.v����a[/�=w��fsI�.������n��w�ن�.9�{8�[h��պ�s�a����W�?�_���GP*��kjg�T��\D��
�,Zճn��,y�xbC{JNL@g�}����Kr�{�,K�;�V�&�E�]+ͽ�G��	�n��S��:�V�F�7���Ӯ �E��Z�����Ԡ�촀����.sz��4��� ��Y��!�';���洄 XK>Ik�svM�DVB�eAx�YO�;/θ�Nv����>Wm����K*���7�4�-鷝�aR���L�ͩ��Pc��z5�w9�x]!�׏(��=��>��é��p�g4����[~�OWg)�Y�ï�;���낈�9���gg�z�t�$���I���<6"��� ۲D����HX��6��}gH�#sL!Es�����s���]A��	����ۃ�Q?���d5�ʈ������}H<�Ń�6��	�~��A6����)��R��� ��v��l �|�t�}:w(��Mח2*Hϙq!e������_�a4�7$k/jt�k��`f�1Ă��O��As_z����v'�6��lbb�*Xj{�O�����ac�'�6�i|����o^������$v~^X�H��� �����B�ʝ˰@iw�u� ��;M~�fF	R�K�׻�02�������q����0I�?0�\?�I��\�N�5��$�l-�?;�"�=��oV�����{��G}W�UG��T��I����ÖR�yQ���`9�K�ҁT�G\B��8/Ľ�~�v�8�Iz����sx~N�?4��!����F9��j6�����>6DE�eJ_�c�{��Vbcp+�rF�������s���|�����f-p#
� ۵�FR�[��^f���,Q҉Cc���k��Q������X�j�$6jƑ2��ȄiT
v���k�:	~�$w�����}�n���6�J�]�E6m����!3+P&s�+�9%㸝��E����ۄ��T�����3��!��ɩ(C�CP��i"��b�=H�w��'�zH�ޡ�k+7�X�e��h�&)��=�B��(���ej�l��� �k�R	�Ά�Vb�p>�y�񤉤4o���!�nِ���?�z�'[TT�{ߍ���)��8���yŪ������^Rs��c$��ӷ<<���V{c]��