XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l���L������m�Nw4�&�o���p|QqV��U]B�B�3bOV�.Hc"Z����R�+�������K��xu�_�o5��}=��n�#ξ�S+���G��v�B�$��[��V�Ǖ�
[�(��m:�U���;z����-S	�́�� �j'�'�7�_�H�~��1��fL*�DK�b�'����,()�������q%?�n�%��
(�ԲeR�3)-GAB$������<��,(�$�xby'e���s��qFV���!�Y/�b(0�}�ܹr8/x�4q�	�#��Z�2̬�e�#�5�A��j~�pS4�N7x�?*��hvI��G�k
Z�3�s��WtG{�������O���;�}�#˻�'陛��5T:i�!�:�����O��-,;]K��e�q���!�s2�w�!12m��=�����j��F.��h�w�9zӃ�#F[DG+��KQ ����J{Z�^+�G�_�F�6�\w�ҟdM l#@�j�Vh�;^�Lo�KT�W�݉�W��>J�n���V�3�ʪ��|�&$�<p���B�E�j̪e5�|V����xN7r[� ��F_���nU-��|	#�Y<e�,��1:�r��
�C������K�`���N!wMx)�s�,�z��\�G��B��sG���쒟�s-����?��v*����׍�.y!4�}�L�v$L;�c�A2�%�:R�����1I�_�?Yu���p��wqV�]��C���n	�e�^
����=�XlxVHYEB    fa00    2470mb��4!1�	��V����3-o�f�Uu3�j�JKz��i��%Tp������ ��7��'$f�a�Z7	�YK�l2��qK�^��)}����oT�Jg*z��=R|�yN��_���*H�<�5��Z0��s`��L���8�E�r-3��0�����:N���ψ1���i0�f� h�|0�#�P4qe�m�yƀ1�7^����
E{�x��-�M�E~���t��s�p%l�+�pۣd\�K��`¨�
��*�ګ�1&�6k�W�0��lΗ���}�S[~�������.Bj%{�C_%�x_D�:&����@�Uh�X7:�I��J }��d~L4��/9	�o�sCd���D���%�w��q����I��Ogc��QT�[�iV��")ǳ�����6l�㚭�vjָ�Ư���;B�W8�l�Y�3���h�#QC�r��^��P��d<��?��'�'y�����Sp��.���g�����yi=�v;�#zo�����)pzQ��|[��s�ְ��}�{���ɳ����ۥ��M�n?��j�Hr����<���X2h�x�D���������Jյꥦ��B
h�@)�:���.�h"8���/��Mfe=���Y)�.�L"ĭC�]i<l�JT�] �֚��%���}!���g[�_Y��i��vH�Dq+z/�?��o�.��y���UF����KQ��w�a���9�;&B�aL-K�h�2q�G�Uo�@�=��Av���hZ�ɮ*x���X�Rel�=$^A:B.K�ɨ�]^��q�����)���tG����J �<�M��`�:[$�C���ـ�zu��gNc���<d��4�ھ���N<��_Q��	c��D�&��e���Ga��)��Y,4Δ}∳�∞��������3�𾸇ٛ�)�|���iՄ>~�c�V��Fȟ���k3_�ȫƫKx���4�.4��J�o�`������2d[�� �F��������=�3�����&��M�l&��nwP&�ǈP�6h�K�/�46�;��Q���ӵ��1���_\L� �Vd-E��S��Q�(�d�Vc�%LX�諉ʁ��4�[�]�#̱����(Sd&�#C������$@���]���7Ƭ*��Ib��-���8ltq?7O��S:�2U�0�f ��<�o��~��n�|]����̯�5,T[[�B:�Z�Qg���1��K�/ߍ}X�P�
�В�h�lΔ-àH���%��"�`φ�Jxd;�0�ZȌ��7;3􊞪��-�d��=N�Y,�o2Ƃcט���~�)��r$4<s]>#K�xFZx�Ug�w�	R�}]a��{��j���T�\�����s�h+���J5��T~���1��󏞈��ͳ���H/���d�f����b#�Э�W�Fl^I6��Dŋ�N�Ʈ�UxO62=[�F�t^[����t:KX��%(�z�a�P3l慏.ڶ�HJbJ��T����q����Gq�V,ǂOid��c���᝶3f�u��y5�ס��eƢ�ƃ���Z�$�m�w(X	s��/���Y$ט�ޯ:]N��m+��W���|�RSk��X�)0��P�f��Y�y����V��ăڽ]K��٬���rz�ڗ�Լ�g�R��B�('��\�g�GΊ8�P��4.r�6�s)��S{��J�O�D�RJ�#k?���!�'�/0��>`I�NҍҠ��٩�at����h�M���������z�;�߰^kU������m��)B��'����C�n��;s	��O8{H'W�]�/SS��BN��y7`½�8DH�.�X,�H@�����7ܓ-���7T����]O���Y4ѴX�,"Cb���	һ��W�+w�$��Aa?l�#v�OO_�U̝,#��E����ν_��.�n9�ˠ�:�����3�;��q��ZzV-éWg��?�p{�/���]e�t�n�Z����']���_rjF~�"�!hV��	��6���M帢*X�`�
C$g�.u,�����H.}�hʙ����G��V@<3�C���rZG��~��O�d8L�V�~�/�Dg���x�������P��)?}�r2(���6�D ����Dgs�[@��/�=+�_�����Ub�c�w)�y��(t��,�� ���G� �JЂ�dwH�#��⯯~�Z�eu������u]Ȼ��ٍ�:
:H�������F#"���{�%�-��ڕ��r?0 ���{��kK7\�q��	^J�h��Ags�ź�&���]H���B.��VEk;�P�_�,i�����f�*�a��?'�9��	�Q:f��K�	��Q�H瀱��:�#�+��K��C��C�rfl�iח���kk.��U��\���U�9'B-��|5k��qnD 4�P��&ǲ��1i:�tS{�ϰ	��G�m�=:����ٯ32}O
���9�X����Y�+&�Y�,����y1�4V�+b֓go�6x!�[�& J��ݧZN� Pۀ�7SS`ǘ�q9�i>�EP?���n��3����>���?�Z���A�7B�>��xX�L�)��S;M�@>?Ri���?{�Ct8�q�T��,Z��2��T���K�)��^����;��� �,���Z������2�F\m������A�j��EMHe����0�zx�1�w�Ֆ��!%� "R}��W���qG��#��.�E���fdDp���r?,�rP_��&��^8���P4C���GЎLs�#j ���p.7.�ف�b��dO�K���Ag�,�Ŝ�Gl��߫ �j�=u��Q�����z`b� �-I�s]j[�O�V��P�&����
�[�KL�P�4.a&��:cR���Quy��:����.�����M �f��٦9�=0,���Y��P��R>�
�,��_Se��>\[��c�����WR�K"�a�Q��/dO3�����+���v�U`�nn�98#0g��%_E�>0o��*L�GAv�A��n
����K�,$�A�VE"�sD���Q�"�J�e�U��
n�C9�"$�>D �.9��\��u"t��n������0s���O��5�����,��c���l&G�^���b����ђ}~��ff./:8W�t�6<��EčdUT�s��}�6i�6�9� /���yȟ�E����O����2�,g�CM9�^1B���2˃��Mn 2��QL��A�c�)&�sx�g�)�#�^�����ʚ_Ok���G{N�z�T%AEh�G�Dck�Op�9r7���'Fb���`T^����ʌ���7�B2�R��vǜ.UC�.1��_G�6��r�u�G˙����r:���.|������EDw�<>�z6eX~��d�{LD���u�0B�5w��0�X�Y9�d�c�h��И$�8xK��V[k�w�J�fq���='�� |�gŕ��v�1M�<%F�.1�Tۍ��M>a��?������a��q�$��j�"7��\��X��o�n�o����C���cA���5gn��&��b�,&+�LtMxD�O,�lٗY�2E�8��(��k���q�h�2V�N��!�A#���r;7�[���qsek7mk��q�2yl}Y������*��3*��]2?�tE�� l\���\�>n��1���)�����������!D-���|G����콞��	b}f�0�*�����t�[�rRS*���3����0I�A�M��k�V���Z�\"���f�~���5X�����y�Nfj��0z$5O��ߑk�����K�g"%�c�;����b+}lg�;4�����V�\X�\xQm�kT�QH�ߝ�������!�O$1Φ�����+ܬb��i{��Ɋ��P�s}~���S�k����h�B�.՟�H3�?�α˞
�`_"��˙����u���/������x�_�uR3f�4g%�_�C����<[ �9�q����%r=U��<.��$�u
�1�/r9�H{��Nq����6��OE����(���05d����uc�_"��P�H9��7%����w�d�e��U���m��|s'|�[ںN�Dd��Z����w7`<r���w������Wɬ�h�)'4�Z���0\ykA�m�]��60���dgS1t<v��|��J���~�}�k�ԋ�����!v��K��P���UQe���8
O*��ܳ����+�ߞ;8�s�,P�(ǈ�G
����o.�<*T#Ӂr4R��kƥ���l�+����v0r��>�7.U[xG�v'y$�k�*�P��w=�]ڿNvM���Դ����W��HcEO��5^��C�)ैL��?7���	���������4R]����2������_���;��U��T�K���^O�����X1WLV�.���K�������7�����(�$ޝ8�i��}���m�c  ���~q(��4�n[Ÿ� \c�Qbh�C�/^��N��K���	�<��b B��3͈�'bv_UI��C2�k>�픆�}�Ռ�6*PW*�|q�|Sa��g��d��A�~%|�������E"djUė��7�}Z���"�|�?Mg1�5NU��(Â���鯗w"	���75��]\&�����~C	���T�Z�dq�Qo�l�\�ɴ�>ѹ����2��.L9�ZN�����Ͽ�0;q#��d�#�	�60:��#^Ş5�RT�_��ϊ��I`�!�WPT�������^_C�\�0��m'���S��j�P���Բjt�{��A��>�Lg�A�f[A^��R�1+�M�5��٣Y<���l��^P�>>m*�0��z;6(��cD�V���SUu�a���?Tz6����~W(p���"�h�51���� &x1�z���\U5!�p���pL4�|��̀���&�^/
[L �/�A)3`{����E�������!u�\Ȉ���\o *_�Up�T��Ȕ i ���Q��*���s��xg8����ޢi&�Լ(a��&�����`�F�y�����3����\V"�>?���)����	�"\zC�D>��Q�Y�n=r���Bk�����i�n� �Q�T� �u�F���eS�K��p��ʖ��M�'�-1sd��Ԍ�i�Ĭ6{�|�[b��߮�3�@�������U�oLZ/Ox�2i_҃{aJ��f�|s<�Ut��z@}�8�m������� R���K>{��<�P/2J*k��2�M�I���NK�rҪ�.d�d%��T�i{�g��������Z�XU��Z�D�6�����Y]�Tp2�t����(��8'D��O�N�"Y(�Z�P���ݬ� �/�"���.`�˿���ٚf��iF/T�aժ�<6�m�}/�������Ԛ���o�� �(]���s�S=Q����0�X�_��w���dey�I>t�3fJ�O��5U2��O��6��e|_@��Fdp�UH=n�~����b�Cx=cW�����$B3(��n�|,�T�}��F��fb|٢ik���/ud�2`����Ŝ,��;�w a�Q`��洒ƌY B�>�u�4$3�2�P+3�:d]��>Vi'lcX��F���N��/Ǳ	]@*�gd�g�dp�y��1��[��~��t��2唣���ޓHh��G�5���~v�����I\q�3�,<I�e�}k�Ѧ����&gxd<o����cZ�%)~���j�:�X�b˟-�T�W�4�
�fk��u�[;+]���]֥!K�������% m%{T���j+VR>�k_Q�_����|�c�*�JT��߲�I�V��n�:���*0<(�__�܇3�;�g뭖�ؓ1"��ys��xS�98Ęğ���V\W��>:��5��N��h$�j����)�@tX�{�����G}�F$_�=���	3�HW_{`g4C���B�A9o���[`u�8��W�PU�5l������j�u�����ˠ�-{�!
E�( ����D��ٌ����$-0$Q�}i�E}�y �A�Z��n>b*57���%��4�� 1uB����ȓ��^|�Wz�i-%��ݠC/�f��S�]*Y��ad�ue$I��0&x�T�ީo0�x��\���Ϭ�:�Ç���j��v��oh�����3��u�5Z�F����.kRߓ ܹ�a��-z�	CQs�a�^ D��N#n#���0��{��)�Q������eaƷ��տ�\�g}��ےC�WM��Q�*o� ֜#�ʁ���՚�D���7�X������2M���%��<�^7,:��O��U��Eb�)���X#^��k�<�@̶��d:ǾVk3��w��Bȁ���o�(��&���ը,'+E}��/6���܀ғnQ��0�Q�!���	��w<�����uRZ�� �1|K�Gڃy�t�����8ʱ�H��ש��h�[*��9B˝"޺�8*�f��g8�A��ir�3�D'�����7��Bz�q�����a���r{�e��2�R,>C>��M���P_^��$v�5E��b� �m����r6=��Y�9��U0��W�4�Ŀ\�(�0c�v�
��&�QЛ���AT%z�+�*���ud�����%��J��n`��nd�M�׀2	P�,L~�Bziʏ���NeG�g��޿F��}~u��|a�x�8J|Ǟ���#n[��D&7PW������O����5��_~����f�Z�@OhT
9�%�"��5pa�Aa�b�괭;{P�;��� �6sWܒ�l��6�đ�륪?��`	�q�U��@y�+̢͸)L��T{W�b>�#�>J�O_F߹e��ucC�2�X�̇~�T�b�o|������C1΁[���1�S�z��ЍOG�W���z�7�+� �x�(���O*Hր^#6�NˏIT⬗�g����#	�b���|��(?j����T�B�\��	D��p1��슺3hrQ?w�1^t�6nh9\�^\��1�&�ʤ\d���fL�r����o��޼�h`���X�����	[�WRM����7`�p��
�U߂��H> 7�Z�ʲ�����s��aJ��	4�7+�����������@V֯��\�W��`�d�Z݅���������Ɔ����{�S$���)'������m[�O���(s;4tc�B1R9�^��𦫬 �����2�e�cM92*e��a+w��_`S����x�2��z���.L4�a����R��j۴s�,�e�����+,��c40���K�~���V�z�WH�Dбs��4
S��1M�Q��K	��s��T]���C�g�����t��~P�p�Fg"G�Z9�]�z-�u�p�5޼%�%��B4�~�]T�J�M;�l�RQY>a���:�-�YU
�:��(�2��B���|�,7J3�.t�xO���{� I��9�({�5�>���!F2t�$��g\�v�_n�w�)���8��%zT�i>��KN�o�qR�'_AYg�Z`� 6}u% �`[�:�*���Mhq�0�s��BA�u%Y�S��(AB��1�+4��K8{��B���O��2`�5a�ɐ<�\=a�k@�1��=�D3a w��^��N��[9_��̲���\ʉp�P��#��{��#�삁�u�`t��B�H��Xo�̤���D7��\g�W_z�i��O�#����zr��9<�m��������\�6�t�ͬN�rx�	�X]7�{�Wv)d/������*���<<V)KT���	���U!����i�y��*sP����q����\6K�"+�B�e�8F.ʬCG�X�邽	�&}z�\�YӲ;�ϔ�b'^<�f����'?��B*���7s�o�����;�OH�Rwe��b�h�ͶI�)c4��� .ά������S��B�/e�r��r�x\�((_�͑�h_�#�l
�n
�yͥ���T7�M.'���hd㑑����>�<Gx�����\D���|S��I�&�Yd���	�h|4.́ >�nFx��G�˜�qX�~N���ٗ|(��W'�G� x{��?Jw�5>k����Y�fa<��c�Ҩ��#IB�T�bzkV�0�S{�=���#��J����J���nq��1؄^c�d;�&���7p$.���� =�{o��LM�h��d�j9nw��������8 B���2��K#2��:��8;���H�SAZgI)J@h��M^�mm��Y��+%�P%w�ӡ.�r��N����ͮ��~>�r����wpG�nb�`N ��-J�W�?�!��f<(�2޹Eo���z7#�U�I OSYU�lOG�x^��SֻḦ�������0���9���9 �Q��i�6F'��6 ��"W3%�l��I�]uW����]�J���z���/�!`�%gn���m/`��<95����A�ZRuܐ$MC?b�C+�J��L��}�d�3�(�F�8�]�?;�$2�d������ʏS�p"||�W���cLX)v�F8� �N 	�1���^�J�g�Esqlb���*}[+ZD$�9�zAn5��m�ۢZh�	�kH����X����S��8.K�^�c-���ؤOB���M�x�w���:���S�q=t��;5m��6�[��U����AP�p���R��L�p���ڛm�ԮrqZ��aˠ���&U�2���c%�V�������.r0�DqMp-�����i+J�������*	���2 �
}����;ǈ�'Sq�ӨJ!B�����
6�rkCƐ��~cB�EW��q���[G���\ru״�DU�K��Hl	L	���AA��]�p8��w�$�4�5e��q���2�J�+14A�q���y��8�#�R����Ǝr���V����+�GX�=V��l�:�M:�",A�	= ɢ[��Α���K�����/���L^��iZB��3�Z����-�����2�+��`��rj�H�r�8S��puO�l��~%�d����/���MTZz%i�g��T�9'}$��5Q�ثv��#Y��HyOH�7[X�j*G �5�F&Vc�j��am�� �0�ĻG�/Gئ��N����@k��L`���|�Kip�C�������	Hj���ť&e/22��^��"+}'A�f"�N�7Wo�}�Z1����u[��OD�^n枧` �8������XlxVHYEB    fa00    1b30#s��PKq���e�7�cs*'*��()2�x�+�y��g��}���n���&�?#�[[*=Lrt����ј�1��aj;〓A��>��8�������|�n�H������"x����!�XG��:$���ף*{J���݀�Q�;?c��~wT�g��%#�<�sr���J����H�bU]�LA���J��Ǣ.�5�&�Y�Fᱡ��Zk%5��Y��j����iΤ���I�9� ~%�%�YΡ���#~�������Ή�Z��ٟY?��x�Svi�J�I�s��1R6��U�B7��Q���$	��O��BU�F����4*�Y�B����7t��ƙ_��㌮<G��+79�M��᥇��/N�25�c�l�m�����Z�Ƅ���ΓU�(��+�vY`y}' �簴4�+�_V�+���������p5���pBd�ҋ��h��V'I��ʭ��+������Z���"xgpJ����@Ɔ/�h�(�d�E��;�_�L��8hpH@k��'|��&fz���xXY�fEb|
��]�ZP��u�זX&$�UJ���dA�{�[)%��6Pzv �-o�~��:�+�c��O�;�_/������ s����4�p��F��D�J�F2GۼU�{�ǎ����sGD\��:C�<?=X����g]�r�7��@���D� �k}���M�B��i�	B-���B�dT���ͮ��fjwP'l�;e�튱��ʺ5�&ޠ8w!f�ߍ�-�$0��b��D��yN1��v\Рa�8^[�]�~URP�#`��N�8�̿X�S���gt�'�\*K	~X�*,�{ogz�Uu�'ά y#_�-R�1���b�ubU��(��ˊG��~o�Y�%��;˰�F�"�E&���ŇB��O�wh��>���y��)��H�L=0�"M/�8s3W�? КJ}ȼ3�
~����ٖ\��l��b2��KM�}qFIR,��>*1,su�(g�)#��m�S��Zޡ��$%Ƒ�*��u�U#��uȞ�R��6�(��p��&��I�8����O�p��r�zk�xuz�����+b�q8�Io�U��|�S皙ARzI�@'f�`�Ί�?%ߴ���Gݬ)ΩtP�E� s�֕o�+�l�6f�l��ǔw�a'|��t�w����'����ͩ˨�����3����[���� �><ak����'<3 !DdJ^�V��Rwq#��3/�d[S=��8!#��_(%�?�b%�7M�A46��h$��X�`R`}�#�}3l��1걚� ����!�g��=Фd�.� �{���j�ϚsK�]W�K�Z�y8��*\��h�fs��{�:�k_b��2bG	��2�s�|�|�=s�j�9H�,��t�}1��LQ�u�?��1�t���j� A�x
�C�¼ۼ��6S gYB�C 4�ҏ�b��Tˎȸ4���qL� /Mb^�;?�N,�"O?�&#��:3�4�H�>�b,�����p��E��+y���|n"�� ވ���X���GN�'Ag��К.^T+�A�-�;2cH��@�G3D��#��dh�H���K��� �����i@��r�{	����q�-ݹ˝� �_����|?$5�!Y��/�\�T.*�z�[����K��	E�e$�Z#!��C�#�|A��V���,�D
T���}R��S�*yAW��"��%�;Q��nE �1�"zY�ڙ����}"�f�V&����N���u�:�-6��Ś~�ߟ���p�CJ7̈́(��\�ߘ2��L�+v��i���e��AR��iƶ�-Tǁ��'�:����,�.�քFB���ɛ_P�F���F��b����+��wEi*�8_���X��_�:=��,_�ڎ-��1�Y��V+���B�3d^5↬ ��-�-�9��?��Um�+�e�y�y���)���VU�%�e�p�k�fSҰd0,�����7��[��2�S�Q#Ɩ�|iQ�;�k���o�i���sȑ}F�/��nc�G`��m�����{���|��ԙY��ݛ+���9��o�T�t��u� �n���qo!�n!�W�b���ףs2i�\�ߧE�bc��kk�r�u�Ǭ��:ep1�*`��Ô"
�:����#<������érypDE~K�#�9����B������VzS�Z�ߢ�n���e�aX�V����p �J���#( �����������Zu���� �K�]�ҍ��P)��K��x赬���>gh��oHo�2q�k>���lǁ����l�t�`�r?���}x�"!)�������/��f��ŧ>�J���9�*���j�v2f���	��
����M�u�J%6Ѐd�z����d�>3��H�GJ���������6A)0O
���tc+%9EP+9l��䓋�"�3��)���D���xݫwke��(��	�rN�����9jloA{0��O� 7L��v�+��gF�Y6�^���5VJ󜽭��䂱��(c�)Gf�7��rd,'N4Dg��宍+-[�*�R�S�b��,J�����@3\2�.r���TI��s(�n�k�+��F±"�
��e����N���q�?��L<�?��TA�r/���O�:�hD5�����tʍ��ʛbDb΢ �yy���l�2яe�}�T�"+I�;�M�s
�L���Ke�*7;Y���a���|+N����n���5�q����w��G{�s�@�t��/<X��^�u_I�H�3��-|;;����}�s �Iq���Ӣ��%O,~=��T�> ������N�����Uƍ+�F]�f�4�����V��_ʸVr�Q��ߐ��H>�l�x;	��`�yy�aH�e����\[O����������nC�}�G���i��?��d��P�`]zt�;��(��Y'�1�c���H�m�9�����*Q�4�2�c���:_[��|V���W��7��h�3���rm����,�9C(�V�j��l�/���2�N��J����0p���� �#�����~[���64_aW���8q�OS��螬��l7pb �nav����<c��������-���Us�XE;��A�H�Z9�}����󂭂���ߙ�ܝ[5�L��`Zg���HoQΣ#��!�n�%�kc�b�h��¯'ZRN�iB��ԫ�3Y~�<Zd�j�u���0tof5��9�}U?\��F�}����t~E+}��^JC�@]|�� ��j�D[(_�NV�d����Y�I�|��H8��?���e��M ����H=;i(* �0�WǕ�9�8#�Q|��"��5��빰aNY{gU,�n0Yؔ/��(��X���|�7��]-��4���ㆣ^yc�����Zi��2��Uƕ��W�x�3W����g�%���+PjTE�E�O>PpY���=gv�:Hٰ@1���"(s{\�z{��[-?�'��=�K��C�U���N�m����񺈈46�C���I���E�2D.�^g��[��Q��^����M�f�B����e��Di���*̨�%vPp�~���y��>j�|��}��y�Ed��?[�{�Z�'��?Le�QyF9\����>X�����t�d��B�EĐY譣|�W(�Ts�O���ȷ�������C����c�R�G%���~�g���,�V	 ���Sλb��h��\�j��ދ�B$�p��iٞ�F� kV���Y,������������Y[��J!dŉk� w[0@�}�3�C�c�"����$�RyrOX�f�}��%-�K-5-fq$f�O=]���A�Ch��B������J���m�_wz���imң�
K�%}KV���o;�%��Z��C��b�����h��cW�5uj��n�|�#�u��^��1eUp3�O���W�u���@o�{�:�-��+,P�ʥ��"�s�f���^�?d�H5��*]��������E
�fV4��f��d|�/�.�����u�bs��Z��7?�sJKfC�҈h��]//rՇ�/���c�XB�%����z��2�����F ���{��+�%G�r�ͯ 0���H�=��UX��h�{�8[�����{��X�Z��WwR��i��4�}�>�4������택T�[?�����!??��%z��goAR�7f��a-o���eX����yަ7�6�7��Oj���Ҵ;��7��;���$n�`�H�4��Ǧ���Fu�V��K�^��b��T���\� �h�l�g���F�E�*�{��d�B^2}������9
��lA�hf�/s��m�*��	����Ђ�5�%9l���mod�/e�ҽ�n���4��{�&~g8��R[)��~�ڱ瞀a�o��$�PoRB�҆ 
NET�H~�{%����t�|'� e�gr��
zo�>�I�`?7rjdBhդ��L�� ���Fu Y�.�K�Gh'�۸�-��uL�~�-�<X��s���2#eSXr���ՠ;�(�2!i�R��#�χ��r����Q����ר�ޒ�J�cP�udb�*�K�Y�ߴf|� g��^���#8�:T���;�t� �7{wI��e+jY�ʭ?�`����I�Y�B��➃�ӵ���~�0�	�l�͍k�~ R�/WQY���ȥe�i��Y|*.��>%�
�c���j�3�.��!Z�����H�4��0�_�X�ų� �����ЏK��,J^��0@�S�|J5�6���QLUQ��e'%D�(�]�t����fk�o{���&8��ԅ/8e>�3�Ƶ�X�Lf%�T�}�n���gTkG+�[0Vu�m+ݐ�/-o�HKxc�;_Km��R9L��h,Ԭ�Xﺃ&;�c���G����������-�0�����UY��UW�,����*'w�;��*�,3��!vZ/	�K���*�<�v�t��C�� wI�Ы`�[M�y�[�q����������8=�޻����)2��i�]	B<�L{�����ȷ��
�t[��U�"Y\JQ�Y���-�0��}��kh���h�ɀҞ	u��)<M�?=b��<77��x��W�]�򠋗��oP�9�4��!=�9J�Q> F�
[Vt��{-k����>�(�9O�s/�h���5r�Ej_��MF��������$�w�mh��S�g�	��Bf'}�?���B ��s��9%9���P0\�k.pC]c9�/��W0&[��I�:%"�ܟ!(�����7+�5�C�P�0��Ѡ[��U�p�M�$�R��\�W�2y���p�Z5x.D�.*:J���0�zG�䍚^-b�P?�-��9���X���>�����]N��R�^�и=�O�azD�b�������	�C�|���s��vƤ�-�"eL�{,�~�n���a�l�*���T������~��"m�reظV�j���p��5j]�Hq�CKٟ�Y��~᮱�kR`��LnX�;�
��B�ފaFAa�Ͽ���܊g�5� ��,?�0!ӟ�t�.��|z���L�M�R�*P_AP�W�B����`�ݤPGN`^W8·�[u��ʸa�E�pRyn���~�)�崛��]`H�߷,�jon�&��<������kBm���I�×�����6���*u�\��IW��;� 8ųTm��Q�!w�ުA�J�l�݃e���I�������������\��Ng�	��ϰ@�=�i��S�%s=ؑ�H�~�B  ա���Y�q�pP\ &�?^M!w[�z���'�=�C
�3�k�
��.��B����H�����6#,i/���ʳ��ďT���+Fd�d�;���7�����`���ǵ�~������٨G��7��&��i���h(l?�!֪:=�gd�K�3��D!_ta��E7�q�VDw����6px"Gx@�P�����{t~,�ƍ	f$M}�5Ao��߱��X�����^4P�^�:_���V&Mr����}�t��Cf���l���C=��I}aX^b7�����R���d���%*gM��6v��_��I���R��?o�Fbz����^�X�0����b��Lh�A��i0���P�M�W,x��T�qInn���GK�l�4�#����O,��i����);x)����j"��w�D���4�@�#{�� t����9I=&�H�Cb`��-��^�#�=�`9�eq@=P��\������5��5˸�1�v[��~��u�{��^.��YT�5���L�.�p!4E9;,�e� �u½�i��أ�e�6H�U�|�Rĉ-�+	�ww������l�'`�-#�'�+y��\� &������=�<���L!Q{]6Hgh��nBp&Y8lK�5W:&w�$�v�<5��]��t;*�=1�%��kF��4HȥR�P�����B+�"�L������,�L���j��D/�Z�&iG��;*�q�V(1��ؾE,��z?�ݡW���־p�NOl��eC�"�0;Z����ȣ�o٧�M]��o��v���0j9�������v�����1\����ȣ�T�5#F�~�~�/ʂn�:F�(+TQ%Ua�ȉ!��9;4$q�(~:���T/J�J\���@i�T'&2�����i	�
wYIE�Y��Q��!cIKCj�'4T�>�pԷ�Tƞ8pi��w����P����u�͓�W�`v�`~k�$7���nB�������S�b��Z=&g��r��9�I�s��2�)Pk+x�XE7�v�O¹��'[}�V�,�(0�t�:���v 2<8,�9H"��ߎ����W��@�'��Y���n9v팲X0�J/��Rk�QE�������L��L�"��|�A�������~ʤq%n�	�XlxVHYEB    fa00    1950�;�"��L��[zʇc���)u�m��s�������K��f{NL2�jf`J-|����S�/*��	7
^�-��e*�`�~�ky)vU��R���W�t��M���h�ъ�en?<�!S�~��L�������4�����d���2�H(��6m��,s)�X��dZ|1?�$�=���t2�K`]�q~Y���PR^x�m4��t�SRe�RH���0���g1+ �������2w���9��?7��y��fsE�z�X��о�_TE3"���^���T��Ir����)�7Ӵ��$Oq@�:��-�!�b�X��;X��T��I���e�f��g�HfD|l]N{���zY��Q���F��I�o���o:�����ȸ�_ч��H��t�	{��0+�9����־�$���\�+Osm����lG��7�+���\�����D��!�J
Q�I���ش���i����D��#�E �C.�D�#��1A� �$V�r���/l�L���4�/[�1����*]&���c(�ϡ،��JE߉Ӊ��_��{�&�����~�Ad��GD�P`r=�F@�ft�O�q���x�n�t���}��␹��Z����|4�Z�~i����g�e�RQ�tW��Ă�O[�[8[����Q�H�$��2�M$K�ϯC���L��h���Q,[�X�d�ױG���q���� A����岗Rb��˂�� ��r��#�l��O+Ƹ[j�)��_�`��lދZW�ۤV�����ص��놪�h��{е=�HCAډGn��{�G��\���u�2����o�4�F$�L�.�4,���i&���*��g�~����~/>��om���} 7t&�aeF����8��K�Q��J�y\���t��?˺�l��������$Q�U�U҃�f�0e�:O�:�Vy s��ga��&�CK���Esy|I���=Jo��jMv�����ϸ���>&`Q�2?p9�,L��1Z��M.�Wj�w�n�+w{v\b��C-F�Ӳ��;2ޤ7�}�9>�U�O/~�2��E_s)&� v�*Y��HI��oˀ�����̳g���Xͻ�X����?��!g���V�+2�#;�o�j;�k�_MU��0V�x�D*CO��H����|XG&��@����?��������6�ށ��q{��X�\�pC�f�u��9��z���D)W�nL��L������z�"����ϣ�Py��T[�g���G���QE���J��W�v}�h<���f�Y�e͐�f�Ҍ�P�/�6�e�'�yl�*@��b'78@U4�a�E}�5%�<Qq�Yy:"�eh�HV|���bZ���&>8L���[m��g?�|,ί��`�n�����R·��$p��,���9Ҙ�(^ȁ�0��T��d��]b��3�u�>*< J:�]�g��9Z. ���C�G�Sjk�V�+����S:�7q3֓p�PP�,���F�tb-7��w��k��(�e^
uV_��_`R�"
K���ox&�|�QS�}�d�!~\�k/<2be����U�#�m�=Q��6��C���2P�AT�Q����՞��d�9bs�Kp�֞������Ύ���ro� ����˽�^�]:�=�{
��ܧ¡4�������?�l�|K�򰮲�����`^��(4��X�u$A� o[��e�X#'����&��L����?d�榡�W`�� ���}@�Gb�	�'uب��y(j�Ǫ!_N7�н�Ӷl=u.ʮ�I�oa�{�?k�k�Ȥq��\���:�y�5�U��i�q��7�^v���:7�J�&�����r��6JDŽ2���Ȋ�3����@Ì�.����ja��`2T�tչ��9�e��5��%�~	�
�8Vl`	�����D�붂��hZ���a雪��x��)2˲�N�w+md&9�����eڴ�����U��-���1���"U�Ӌ%��S��u�̱�yh1������2*ޖ88�0s���������A8��x;��*��y� �O�u?�eQ���Bќ[���N�k#��Va��م-�R���b0gx���P�������UVsZ"�E�s�9[��߷�-&#�p�z���?�_1��ۈ_Z�*� i�ۮ�aFyM2��:tB�	s��f��n����v�R��	?V�@4*Pu����L�jՓ�����Z��������������4��M����#U)Q��X@/������f {�xW�8_�B���*�1�ޒ����tJ�(����+߂#�p+'�i�f&�V`^t�Z�j!�ɑ�;`� ��UB����J�k������,����[���P��yǲ@����u��D�����CV���|�a���������6��oW�"�e�"��J�}��AO�Sk9���K��kḀ�z��d�E����?+1e"�$��0qi�ݬ�j���5��Ku�]����-��E֞S����cq��K�Iiˡ�g�h���#®��������[�H:���ȯۖ��[�ͻ���jd�����8pG���(�8�o'oG�=���3�}�
�e/� ��K#м���^���6� O�pV�x��a�㤪v�O��^�REǒ\׵�����W�'��և��MA(���s�L^�v�U���?��g��.xgP뉓�F�ʾS�^��D�4�%��H*l��4�;�ChPqp�xH�3��Ӣ�U^�sE$�Ҏ�2���69��p#�7��SD:xQ� ��*�nTͻI"�?�A̧����HmGШ�2V|hǽj�2̵5����l�D
��n��+��b���\GyK3t`_<y��K���3gr$�͟��$bh��-\�;WxWj��7�v��II�`)Q��+��,�E�oLk��<��X_�-���K�� �t��j�I{� �	���
c�#�[�u�<�_J���t���d�]����Z&��Z�#}�\�ެZ��)��b��\�I�?E�Q�x�Kڱ7ˢ�xԟ� <w!��n���7Y�N�;J��Y;���\�i ��N6�r�̽�AK|�9#�bZ��캞K^^w��Dj����:cM�Wy� ����kܻ��0-�K4k�J|㸯@�s��kN�k�� ۸�GqdY��i�JÇHjF[v� #�2���<(�/� ���SH@p��������Ѧ4��p�^�Za�H�4�����37�R*�|7�S�@��S�����\=�U��w*ܠ���3���ƭ��/ݗ/e�R[�m��$��loN*̌�3pij��
K_�����pv҅6s�o0	2�׭�3঵�v��c�����=B�L��Pu2#w���?M�sm#�W�|�c{g���{ɴ����h�������
��JDf�f��Z��-Ϩ%�]F��jK�ԝN�]OJ �n!�K��l�P���aҟ/ܖD3��Ac5�+�p彫o2�=iY���g�����&��yf&V�Y�X�i��$w�w�s�w���^���x�O6�n����8ׁm���Q�ݜA�,��(Suo���
F�b%־X2���~6h ܍$��D�+�����j��b|��Ir�xP\]]�^{�w7.)���u�%�� GaO�F�?�9P��Ζ���s�So�Ύx���L~Y�zCw���9�K�Lݨm�	E�VUտL_���N��z?�*����<t����(��@Y�!@�s�A_i����-�Iva�����Su�6��5�M�`9�t'���}�/-�s������g���S������t[���9B3*UG)h7XW���0)�+̏T�yY��c~�m��Ĕa{�C+�J=T�(��ÿY�X�e?.��;f�x�%���\(����L-s�1i�"����2}=4�K�bD��K��>� @�\��Ot�S��h�t�Dk�����nE�FC����#�m�b��M$储�S�.�Gj�"��p�h��Ua�>�']�<��-F��z+9h�9��F�
/�O.�w[59�q�QM��E��e�%���w]�7/�$����D��x7=�`s�[���HY�,�c_����%�퀥B~K���-�s������Q�w��F�Kǆ�U�suՒ�1����k�L�#O�@lX�\�C(:���v����+I�F��`���ש�5��l��4O����C,��MS�����A9�V��⨍���^��-�DQ���Q1��ptR��l�K�3o�TS��xv7P����������N������X(���A��B��\O+Q����`������{��/o��f���'�g�{����g�������1|�ٺٲ�]W��� ����k��նB�4� ������Wӥ�@X�G�8_��>{S)	1�|��Xٷ�u��)�rk�I%%����k�#����д|�B��,ou3����5[M���|��n���=�D��=,Ňh��e�����Hj������F�w4�����4.�(k�]1yk?���`��F��G�]-��&�b�M�
�{���+����2��-D�����ux]WZ�Ө/$��Fk`��*ND6����[�VL\?{@��h���_\�����y��p�������|�/	?)���mU.�w
:��p�(��^��y�L�3F�w��D`�܌��)�r^K0��Ğ�#n^h�p�q�0�<�i�u�O���\��@0�R�M����"�0As��1 t�Zj�-֣f�1��q>@���ۨs�ŭ"�mr,_��B�|QOB��G�ˉ�z���t�I(�BSގ��*�sdi�Chv����uI@�(�:0qh�/�1;�.���6��Q<��"_�T�wZN�rH���9��w�0��s�ȕ^F]��&'��Dt2�1�	��n�>HL�wj$<9$i L�F�1z�
9��q`�U+�.��E����.*d@�55�s&�1Mo�"W�|�C�W�V����(j�ũFu�,-�c�/B�)�;}=�(�)$��.6��=t�0�^ØY,j�q�S	�%5X'�=��A<��A�!w�0TI��W���į�4ʪ0�7�����O|�{�{����� 9��T���ݳet���`Y�/�;���~�8���z��G �k���o�V�X�'E5:����M:�[Ƥ�Om4�0�{>L�� j���ޏ�K]��#����e�:�0}�GiU�uyv5�l�
ei^dSy5�838�����y�
i�N�a\Dgj�����	ɑ�`ۭ�1����-��A�{o��pa�X�F�N���s���ؗ��q�:�dd���}����cd�=�0���b�w��֡����\�-8~wu3��\9,�R��̮b�T�'�5R��σ��a�c�B����{|�P�-���ĕ�E2���(�:�~�`�ΐ�Z{ma���'_G�״�c3�Q3�ZmhѸm�R��YR@�h%�����^�ǲ��nd�P�Ǉ�K��v�>��ԥ{�����N����j|w*��:�8���PtF�{��v �Mb�)�Tt�ګ_�<A��@Ɇ�6Ҋ6։@����A�x�1�1�(��r�s���u*9r3��׊dǷ�Z8���B����1��m�N]�Ci��x����*7�� ����a�_��'a�Dj������K���ͥ�ވ7�gP���Z�WY
�p�&��ߐP@�Q"5Sŗ�-H%�2p>�Y�ˢx�]}������˫hL���g�P��H��k)�3���Z$i֕۲�	H����a��+�����]	Y�;��|w����N�q�:\X�9㶩{�c7��-h�^џ?�ࡨxW�����hS����4є�P�K��i ��bcڅ��m�`��W�C��2�R�` ݜ����։@%�&G?7i�B���Pf������2�4�h�� {�E��݌	�j��f���ڍ�Ϫ��I=����.�!�h�������)*q���'�M#���f���颫X�9hs�N����7QRY""��&�G<`dGr�j����f/k�/ڔ;����P�0Z�}3��3�Eх0/-S/0��M]Ity�3���v�K�x}2o���G��ő��!Z����K��;hJ-���53�h�E�I m����4���Y���s{�p(�w�&#�Ō��O[ʷ�Z��L���0¢�3�DNDh�:Uo�ֶ�XG�"�0楱ͯ��� �ʡ�/��Y̿��-��L7�����i��?+3�ы�Q�L%>"�ϑ����P"�j��\gۘ��C�g���ܾ�qj�e?��x))�RNKӋՠ�C ���*-V$���V#�9S�/��k�ʰ��V���8��W�@<�0��R��-x�a��XlxVHYEB    4f27     d40m��a�*pФ�|YO֊,�&˘6��Eo�V�{�BL{K$��[��㟹�A5�e�p@��K�9�b�"x��gkD���X��Z�<����xn�g�(��9��9��b�}��l�A��޾y/��J(�1I�8�M�P^1�K�J}��lT �<T�5��oE1���<�t�0�w]HCf�}[E6�M��ѽ�����m�����B68�0�T�)�aN��\ �<��^ja�ϡ���&���\�h9o�mբg�@�M�=�p,�0q!w���Ze����@���|��a�%���/L�s��_*Q_>�r\Ȝ`7F#��B6j�ZH�_��^d�|�� �E ��"1a�Rx%or�`�f��Gݨ��$*^'8J��V���O�Rqe	��S�osR��@���Q-W��eG*����Z*�:1ix-�]`�_�g�U.w}b�0�o����+����?�'�[�5Ţ�A�0�3vn������m�N����EQ"*�(��.��z7�	�l�f�}���k3�8I�k҅,y�$�h������ND��BR�Z8�Rh�2�n8]�#�y4@����5���,�����ң�3����ggٞ�Qm�
�դݰ˼@vlFq!{�7�ʺ��Ym9���ri�-��\浘����w�J
C�yxk��Ό���~(7�A��|�ƶ� 9$�ƺ�$j:i�Ek�R�"LJ1c��z7��`㟑h9������f1"�����є��|��w��Fa�\�}���~P�yM�.��Pf8=>)�G*���0����@�9)�V=����6A�� v��y���Xm���m�N�ȍ{���u30��%����9$�Uy��&�tOk3�C�n<�6؃��[�����I�����`��Õ��7Y�wS�(G�Q(B)����L�S;;?�?`��� ���s�Jk�:��!�~?_G$
��o"��%�j�X8��2R�R�r	�k�9œ�W��N��a�Y%n�QT��RS�$�a�������:�����QE�5_�#<N&�6A����	��@���|��j�l��7�W8�N�{��Jg`o�������<�?*��[�O���{���l�;��L�O��$>ƺ�]f81c��VN�A̚!�B�����[�\W'a��t�cJ��\U�zE��p���8�w��ņ��o�]=.F#}�s3��_�� �m|�U��WPf�c�lvE��/��w�T��j�\�����=h�d@fL�Rt���_�䟑���g5�x��<Ϙ���Y����^m���8՗�A�9�lm�/pJe��={X���G�n~�G.��yH��-��}u���-����Prǝ�~�.~̩$����հ4��*�#������*T
����J߮P�j4R�3H��kG[W��ѷ��Q�	[�� �*��iA��&t]T5"�_G	^O
�wu�\1yt�{�c�c�W�ʫN
�%4X�4Hi����b@Z��Ǆ-׃�Pt��E�Y��r�ĭK�n9�(r��0q��aጴ�c�*E{�P�Ѥ_�����P���4Xq� �_�Ւ����/L�� uB�+���g��"��n�	��[�v��\�F������6�Ӗ��Bؽ$�+@�$�k~&v_XȮ�l���2��@��]>�?RM�u�sA��܆�4V~c֠�[��eԨ��[��/g^r�P|�k�Mm˯����y��� A?F���7�
p����M:���,p�N�����w ?��-R�aq���3N�rRH��7�ňrU�&$�v���)��&�9�UUL�?�⢦O�B�& ꣢뼭�Ӛ�o��(��*���A�s�dǲ��C+56��o2��Q��#ö�W-B3I�ʺ�MY���`}�@�|z�n^�]'z�����]������gk�ً�9�Ux�d��B����~�Of�LlΜb�!���IdͲ�r�[��K �`�<ʍ1��)(����RԵs�TJ$0ҌFU�*�Nu�0H�b�����cs���t2�TJ��U0к~�rGT�����_X�S��B[��Gq�h����Wy�ڂ�+%�GOHcu�u�F,�]��r�:�vĆɐ�p�_�8pdo9����ҿ`a]��rI`�Y�m�K��_�
�ЁuvW�W��� @�_ĺWQN*�!��d����O�д7�n��4��(�,xV/�p��k��s��z��T��|����"�P/]a������$Ζ%Ϟ2�Zq���=�\A��`�k&u�#�4�x,X�]���<�N��"[�+�\'�[�[2�w0�,LU�"�;��}w���a��0���=��9ҫƽ!��>	 �΁����2KІ�;����ͽ1KIJXS����]�`v����\:ZY[���t񫎼�}���
<���18<���QxG��5��J�D]�ia"�Ŕ���aL\��iG���-�s��l��j�P�%�m8�a?�z�T�1O� $��͆�i)4��G^�ٿ�rG@����_4���q���xʲ��i`H�d{�$#$0�:K<Р�������j-R�8�b��˂urp]�hQe�E������4s�����
�>���եD��Sp�M-cV} ��ٽ0�*:��'E���U��t��0�'�ּ��Rnl�Mn����&lK�V��ᾘ�٬��3-��>q�"_�����8��&QȤW�ٽ��^�j�]��gJ�M�s;UV\�[���$VX��0�+Z܈V�?d����
)J
�����ܲ��-M�����#��|Z�����y)�@�r�v85�X�d�~*�}z�~4�=gǗ����y�'����C��4��I�V�7TT(Y�:���LP�և�ԋ-mM�?�W����?֔Ps����+��/��A���]&28V�R�"����''�=�-����U�S�����L���V��Ͽ_Ͽ���I�D#�L6�6��`���&���5�&�����6� �&Q�+#H6�bk"B��p-ҝE�#TbH�#*���r�/��5���z����eu�U��#mI��b��c� Yُu%,�tsF�7�O� ����AWۏɐ�-&�N� Rz������d�)�s��RZ���L�M�r_��(Ho��0|+f4��Zh�LB�sPz��R2rkmUֲ�/�y[�	ڏuM�_+�13�R��)~Jy` ~�k<�3z_�;�m_}��38n����~_ErQ3, ir4e���w_�}+�R��A
�V!뉌6�m�7�Z���ѽ7ڴ�����j�;k�ֈ��>�r��E2�c����̘:h��ۖ )�*SaLv*��RC��I\gcO<�^�%H'�