XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AL�n�0D������\V~���+ݎA����!�{ZS`1>�9.#0�j� F\��$�������VKon:�VĽ�,Ӝw9 }�\B�j��t�[;�U�#Ĩ�s��p��F���Ǐ�P}�9X�jBM����[����9��yA�{_"d��$��z� $�k4� mW^����R#ϱ*�~⎛�Ex��UD��T�r9n��-|�=7BQ���5ß@�GƚPƘ�7xj��e����C� ���rӏ�A.'md�V��j9��U�`�f�F��'��w�Х}�
Dze�ʍ�R��~'��i�ڀ���bt���Ux�Z%zcU|�j�7dk͎GX^����k�Y5���3��ו�Z ��$��w�>I�֑຀�}�U����a̶��M��n�7�+O#^�Z�� Z-I�4o	��T֧9�ݣ�p�>r�X�:"�­�=Yidm�J��"�n�� �#�n���	�k��P��ڢ��\���D}��2��m2i���u�:u�T��Ӆ��D��[������+�h~6BOES�sm%�Jm����?�(0O��m����>��NDr����7���}1��[Eܘ�F�H��!�x��IJ*�6�sl�3�V.X�p |�bӥ)	�G!U�l��Fh�K�i�<�� ��f��oA%dxe��:�B�iz^�[ ŕ| >���u7K�沓n�2����9Nȼ�r��淒�Qm��X�>~U����u/�X��4��uΥ����YL�Y8���XlxVHYEB    c3e8    1d20/J��T�*�]�G�{�^�{r�S���<]4�������UY�`�(�?�9$�e�j�@u
�\���<��C}��4ډ<Zo��~tkoJ_yA�{�r�v�ҥ�=B��ZI4Yz���T܃�<�d�e�΂��$��VUC3����3���i��a.�Fm��9�����@�m�
�������JU�u����2��a���B�ג&S�Y�(��>�.=F�~��R��$N��wIH�<Q7[x^v���(�I,R���h�¨xr����>(}���l~�̰�Ѥ�@��;�X����r.>�Q�%��6�n�/�e�~:�lGr?�H`�����Z+^xa�"��V��3��2���H2��xN��S� ��E�s��po?�31�E�4u��(���.K�X��ތ�p�j�I`˨�����}*�24��$\��T�&��q�:�(J~��ǊWE�7G��5��:Ew=�nf�l�j��M���okoHP��ˎ�i�5�>�b���7b�=�����C��S������3Q����h�K�jG���:�H�;��bA��������1םk'$�J�R�G<L92J3�G�f�,}�M��0m=|���k,Z��f���v{�T�8��H��'-B�C���+tJ-��.�
�w���<i�O���m�^{6QA�F�8dоB�t���;9Uy�'�p+6=�~�7+O@aBt��I�O��[��tW�t �����?^���j��%Ԗ���'�PjJ�_K����c(O?��)��`��	�����I�^ª�qY��DIͮ��`�X�QI��3��)
J�O�s�g����F>�8��	@V*L>:'��!��= $���`��d�n�!�V?sa1ӣ ��n��S�g��^����7o��(%��?��뿋�C�#(�������x��E���@��7 l9p"����f�-��:Am�������<}X_g	���`]7��H�������D��.KF���/Dt�cF�%Cp@<�1d͉������LR7��6ؒ#� ��4[�ƫqr���b�A��|�bmNw��>�K��H�����yn�86)�R�?�����T�]	�-e%TB�<���U�DQ�� G~�ԓ wRֿ�fwD�oJlw#�QMf�z�7�����K=T3�	�|z�n[rn���;a�2��O����A?�D�.x�]p7܀����6n�ߟ�H�Xw�o�ha_�T�~��n'�+!R����$1���ٿd��k���M07���σ�Յ�3L���nJ3�((q��.�8�,-A<XR� YWo�tIdGe���k9��,�-�U��y���d�#$Y��.��(��u�Cv�(�Ԋ��KЗ��|'�{�K����.\�4�Ж��UH��"-cJ���֠�ׂu���3�@�~?���kq肠����߾6�-T}o�z����c�_�is���k��DBP��y�@f[c-��ȑ�Y�M�,(�����gz� �n�D���:�{��yuOl�8����7hV����P!�PVU�9���G�&n0(�S.���y����[��o]��<t�[	|��:p���|Ү9s*$ ���*�$�JJ�{օ��'�&�b�u퐅Td�R��:b���X2�L��9��K��(�N��T�f�7Qp6xH$vD�?:��Zo��c|�VimIg>�������	� �����ڃ�R������EX���]f�T�b���<� nޞ��Hd��*I�׾�E8�����Q��C00�?P"<�E2 6=�Ґ��n����g�_��O��A&�ՔYwq�W�K���-i���W�Me��'���I��_����T�wY�8f�]ۉ���ݙ���`�s�n}Jy7��|]�K!te�S%"w���|df�<�����hz�ke��	�<7�v·�Kb��5;`4/�n�Fr�W6�6��]�%�.����t��/C����
�1�8�[�����	��/��@�@��lT���sW2C�n���u�u��'�UI��1c�ndF�n���0ݓ��ZT~v�:7�Lf��9�ԭ��F�^�[0�G�����������g��*܇�,T?Ʈs�2���A��5������-	��e2��M�j�ZGtC�+�Y�w:����`�T:t��C'���YP<d(}i
v�A�8�P��� :K��o�T֤P��i��F4��<�]Z�/F�[y|oC+mjD����`S�#�5�βOY��9���O_*!���Ω8m=h	��}-}ڍd�QSP���dq`1TFY%Q��7�y��E�wa@�3�A�� '/��4$wNjwqXA�e}}Ԧ��Eg�f���29�H�9�:�ߤ@�$.�j!UZ 6xy׏.�s��n��`h�Mܲ'��v4|\����2A�4r~9��>���E��C<^1�[�2(��6��8{n��8��O��ˇ�t���!�S��*$�%h8'������l���.0{��P�r���EL�����ɽ`��^����$��`n*���F��u���$o�;Ì����vm�^-15K��u;��x�e�z@!���!GG�ᥪdI`���L�5o"'Q�hm���q\��|��jU@�ph, �>��_�%sF��.��rw�mϮ�s5�>�R���WP[w�r ��-�z���F7<��V����NGS���(J\��yD߮��Q:[��o2&�q��kx)t�?�y|(��_����� $�e�_ф�ʷy�����_��М��dױ}c��z�B�+0����/��'�� B�2 T�\3�	I�/��#̙h�7rp��i��rfw��B��5s�Lp�E$&X�sn�7^���)��p�%v4����ˤE�f�2�m;��Y[�^� �D��
��l���^n�`ǂ^����j^�7r���U��� ��/MVL�ܺ݌����Pn�sk�c��*���l+S��/�/�0-��&ubT!F����"꣌=Dth����:��Ix���7XN�=E���g��E[�P�z*���|����I���E���XB�bZ�T
.����9���X���e�:M�U�R����ܠ1WJ93��.��{3 �<�&m>]���	qr�y�/-��WCسy
�'~b\�5E�� N7��y�D�ަUrC; vf��'h���I�:3��TIY`�!��Jx&��z�X�k�9>]�y�'j��g�k�X��!)�[���e��6)�s��}"V��0u&�U+{<]+�!�bٱD�!
��)�V�P&|��d-ƍ-~�Lf`g)"t����,F�i�Ֆ8�V��e�`y�:񿐍`���q��_)~�jE[�6��v>B��k��-1�؄nQ���h������vM�.�����Ew��W�1���ah��F/����[����D �m���0�!Ԇ�@uH�عo|��=M�3Wt��Dq�\f�=؍����P�~�����z�f�r+�������>]�s���)�L����Y�H�ї ������nF�%� PP��W����E6�D`�1��Y6c��>���������/~a��k����f��8Ó��.�\��f7��~ʟr���pm?y�/��j��n���+~:�P�?A�J�!�=��`�|����\�C��?�`�PE�\��}r �R.�Z�a�?>�A+�B�x������	��)oքL����H��ʪT�i���N�]ڧ����;E|��\���_����0k1[���
C����8SR �ɼ�X�8�},�³,��|?9���Pa��*Q����f�&�r�h�X����*�4�z���)�l|����w�V�J�����,|�{Ŧ����KrM�?���^�\n˴�����b�j�{�NRtñ�\�|��rpd[P��lۋV.�����K�֖��%3�+ahD�ىt��^*,ἦ�`N�Gɨ��R!@���L��y��毹��<˺���QPR&���?b��y��O�:I�L׬<���4��I��}<uw�<�J�o[p�,E��Ks��I��Ḽ@�J�Jޜ���YF7rD�E��ˏ'h5������Ml#�"��i���4������3!Av�
���
�
��`���D�N��xz!�(�s�y�J)NG�H�^/�n�P�W`��|٬�S�dc/v��^C+�3CC��_©6�1�3z��/w8���)1�J
G�&�Q?]��-b���Il�Irw���)^��oq����0-�I0�v�x�_}�cCU��#�i��1�����޶�?.\��z�2y��'�hl�BL�DC�����" �T\ѕ�|�܋�J����l��	�"8>\���Ri8>�Xw�%`��gGk�W��'o�4�]��/��D��E�X+Q���ˈ5b�Ag�Dޑ�OIH�򳇸���'Fݶ�"���e_���#���#�ANk���ۅ�`�55�L�x�������\�~�qA���|�;�;گ-�@�V�eC^|ks�\Mt�����<mcSo��+� �����o����N\-U�~Y�G��=�b%#�Z��m��gޔ%n5�K{��ȕ�q��2��x[��(.���������<���Qxm�	R�K���K1�ׅ�<
+mO�_�!Q�!�����A�*�X7���D	zH�և� �>�/
{د݅��$�N������'��+Ñք��D�q�x_9��i*��
�g�q���n�R�~�ÄV�m�FQ����d|%�o����@�a~GO�
���M���7»c�4x�r��fk���&��K�f�|�ڿ��(�������}�hZ���O�U�h���1��g&� j��QK>0� aǘ��.��>H0�����IF�T�e��/r"ư���>d\����.֝��H�r�F��θ�4�R,X`��-�#Jr��ІT�fxc�:4F3�"��3�!�˚��kήtg��s{e����E���C�ˮl/����d����F�,�"0F�4MR4���W��䭲S�E��_�j�9c-�]�v^�yM��Y�3�M����=�Sք���΁G9u�{Xc jkFb@��Mut��Tx�e{ՙF����%ʕ�c���(��*��i���� �ہ;����"��LK0A��pw�%�f�56\��R������ǩLb�g�#��$�N�p��(_���<_p4�Ĕ�Mb�Ӌ��D�W�rLhy��.�Q����_5�l�%-=���Eo1}����'D�&�w2K+ٵF$4r��@�^n�$�8v�d�����1�������M^_��9����N�U���K�Mj`�,��Yg��?h3e������n^`@�%���2��r}q��4�$	Kݪ� �v`Xa<�O�u�f�e@W��l8��mS�T��,��0����szbv*DBM =�����*�0����C�tGz`���l����(�[<�Ӹ*=��K�B�^ Z̘# ˓(�.��h�k@��s�⚀Q��G(6G�e[��}u�]������_�}$%���#
r���N��N�{����a�@�����WƑ�Q
۳۫M,����b�|��z�dj^B<"yU@9^$���I{8̲`
SlD�+�q8b�^��N]*p���
h߃g��k��rQ��u`�b�s�&�V�)U6a�B���%��=~��`�h-O�g4c������v��f��g�Xu�t�l)?[�Z��t��ff��U�#|*�3�~�Kc'�/_�)�XW�3���G��t�'�\��4� ��"q�ui�M�䅊�9F�J�����A�9��)�'����;(~�h�4pd���xf�{�"5l�C����pTp%�
<½�葇*?���}��A�4۩�Lb�\�C�Ӭ�9�y\����ٶC��8�O�l�j�@(諚��f~JT�U����Ԏ�l��5>7.tm]�c�<h"�-�#�uj��ʽ�ܤ�t$L\o�U�3o��E��ṣF��r�ɘ�L�cr;�*��d�[����O>�DLﭒ���q�i?S=3L���-�1E�.$�]$a��o�@��K�0$(�U!|��O�U�����I_������(�J2��e�����_<}?+m�\�0T����Y�A���:�Vyp�4���mؠ�RbT�ZYC|��8�c��H�Y�M�
��8����JE�_�ߢ6�է�
FHH�qE;f�7��:�j0@�bF~���`b��l
e��&:��x�B��
�� ���`9ٷ͸*L})@��4�l��J������S�o�TLϴ�����",S��vqn�h���W�<��H�U��C�@4�	s?��Ĳ8�G�߂^9)� ܘ���]�d-KW�o���4�x~�?�ᆦ� ��M�n9?���u�C�K�u;��?q���{�v]qQ��c��=^$2�t�}����F����,�@Lp�����<~-o�Eo�Q��3�'��B��ՙ�8�9S%�6�*!�>T�q#����Q�ƥ���/^ǊI�zY��^�%e����x�-�G�A�W���o�{.�M�X�C���Zm��k��,�&�w��c����i�����]|x�J:�+~��9�������C�cܞm	�^���4�B����t�K}���ѿ۬�ƕF�I��r���J���um�`��'��jA���|��*�I?�lF�c�me�ñ���jN�?>O���p8��d��GF]3���xU��	�,0L�=a��C�s�8���^�ۆl����L^IQ	��D�~5�pcS�EnI��Ͻ�k����ƌ�gV��7��@Q1�a�g�{�'�����6U��4�ޥ^���T�:�:� �A@��v`j�����e�LO�g�E�z�!.�@�-J͐��)j�Y���2b[��S������"ˁV����O�魂���?	9J�q��I:
�8dӓ'��ރ�g*�ψ��Ѩo݋�~p��VV�V��o�d^2���قvus�%�oMgA�`<�UA5忀y�ߙ@�i9�VFS�8-��r������0yX������0eި��^q�Do��Vĉ�h�������,��-Uh?:�����zC�'��]�0F]��BuF�q��ϒ4�2��$���)lc�V���@ߕ���{ݘ����R���!f��� ���Y���ؐ�����̶��,0�$�Ź�3Q=�!�w)�5H#�@,������0W�L���uIJ�YꇉU����['���UW��&�+�mAB�z������Օ�A<��SAReKSS�^�3���:"����Ns��6k^��A.�� z�ꥊ�{#��H��by&%�(����0זS[w��̨�L$H0��{V7���$3['�x�v�=�G{T��q��2X`��