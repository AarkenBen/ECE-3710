XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Of����"�qV;�p��[���޾�@e�~�.n2u{`�S���|@~rOI<������~͠2|�
:�E�T���C���S��2a�I�-3eǁ/i�\���L�M&�����
�c�ʗ����d��T@�j ����xZP�'-�^8�:�!�nE0�:��\>̟���tڌI*!����g����i�.�OW��b��(�Z�Y�o�Y���
C�X�F8W��aG��W�B�;���t<�!�B�#�&I-n
�Li��)���R��x�E���:^��o���:F�s"ځB�K4�@�u��� �yL#˲���+�1|ٺ������c&o�����6�e�␙��9n�������a��Fs}�y��D���ЀKu�o�^ֹh �;��μ_"f7�,BpK��1� �`a:b&�=�|�isG#��;��س_���Z���� }
�\�����v����?mr�\����!8 ��0n�s��t-��v�����D���� ��D׭��/��s@׊��4;�ێ���c�R�����OεF�7���$�vت}u�|T��� �֫�e��
�褱�}-G�)�%x>�G����I(�t�p�+���$��h��D��Ca���Ҵ+6��(���s?���&Q�_r�|��qC>���d��R{o��I�A�Л��J�6�g��ϴ�17&�2�������_*/3�WV~�Tk67�|��$������'Sa|1O�)�S�T�=%XlxVHYEB    7744    1780 �Yz�ޡ���l�����
hʤ�����3�r#!Ш�F�
�f\�oS�K�87���=(�]������,T�)��69�q0����?d�"{�a���l�gP���09�e
6B���ۨ��3r�<�bdm��<�._~J1,K�hW�fV��N��|��)�4�g�.�j�_�v|������v1,3�YbХT�gk�y��dJ�k�m�d>��R��BP2���\i���9�׽���Bʍ2.�rAƏ�]�;�=�`�!����B������rHl�eHޕ��:II�'��Pz��$����B	O�j�l���҉�,N
��:�2�n$,���+����9�}�L��.�2�yX+ʡ�`.[����j߽���0P�$^֝X�eg���wyx�Q�z��d+���?�n\�iw�ke���mU�m��c�x�E����M�=�Z}�����-�d���q@�����1́!�h�!�r��z꞊�t�v����b�ҹ��?�Hk����p����#K{�i��/�O6�ze��6���6���3z��~ę��#i�߼��5]�AP�([���EV���L�=u#�1�Z4�����4&% 3�_,���i�,ȶ���X胗K�j�?�Z񮍲R$8:�8S�:Ɓ�;�Cr�N~�[cF3�V�֧�.S�/a�15^Z8Tp�bO���s�eɽ�8���������y���E�6;R;�6�F墫����;�� �Q�c���ꗂ��J;L���#ByjC����/�,2�ڼ��عۣ�S	��R���r�˃��ݐG�8]ȵ5W�7��y����jć<��.�����ͫYi��I�#�W��ԑ�W��W�V��&QZ+8�oᑗ�|�?*a���'>�!Ӳl�ϟ:c�m����%|!�G�H�����k�O�q�3����\%T��71��F "��x�$������޳%�H��B������?
Zy���	�}�d����2���y,�y�q�a:>�[�Xw�����A�L��=��q��ů	=F=B��	�y��ȼ�
[9���7�ێ�lD>c�4A�둽�"VZ�߬�-�'���z���ȫ3�/����{:�a�Df�Q��%��H��L�;s�=��?׈"wv�zQ
�N{��JH}p�DP�t�� u�~��G��R�R�u�YyUo��7�P${��0	�R�u�v��{����f�9?e��X�G��d��}�/��s� ogcn��+K�Ӷyv�I߅ZY4<#����z�'|
�{�O�.��:tX��n?x!�r��!E�wMG��k�*�Rv0���K�@��ŭn�k���%�@J����75�sSm���w�>RW�ei{�<U�"46agY��7@�Y�Z����RA�47zH2y�|��XĮ�ZE�ȌŬC���T��"�h�aڹ��Ǟ��5<N�[|T´v-�Ȭ��t(��������7�������w�����S�\��PD!I��|"�"�PW��%��o�<�M5�C�Vx���Gu�~���Վ����=֪�gV��0G3U��^%�
�{o���`���L-
�2ХVm��e �U�kk{%�e�ԕ��P������p�B/�X�H�kd�����;���<�C�+�5��X��h$5��o�����&��a��C"�F��mա~`�VY�t�7�hҜdM��ݖ����y�&����^ʯo�`��B�����	��
j����#�������1��F�%uyI���ьŘ�_w�!��qk�a��M HT8g��a��݅�r�-:|�D�HRxȬS�-*�=3."۫��B��(���|W���h�-�W�uHlF�.����s�6���Ks���,*0���gR}͂���z�����&��d�bX��E׃���Kq�R�f�Ӱ��)�њ�E��@-�E~���N��q�Z��h�h>���Z��-��/����!�Uv=G��&;{I�M�I�/�+�y�[��?lޅ9�4�����`�_X�j5�'?����Ap�p��	B9\��
��@!�_�|�kG�lRe�f��	�� 1��Id�~��o�։�a����W��)�r�#t���R���uV=��jS��� ����(|G`�~�hQ���J䂲Ż����԰2���pIV�30&�u�< ץ���� �  =�M�ձ����u@��r+7�������D�C��Ӕ٧�F֝?��0*�e���6��LM�L��"M&�k�#lG���CmU�Sؒh�Z�c�J4�Q�i˖���e��C�^l���業�o+I�M#�����m~��){mMg����Q�9���_�<���
������u�aЁ�#��[չ[�W��X> ���#���H�^X�(���Q�;a���,���š����S�He��K�t�+�ry)G�Ds�I�F��Av���ϭ
6'����-vnɄ��P��u�X@�\�|�b�N(���7w��S,�U��ݜ��]�+�XJ�\���0*�R����`�d�v�?�ޗ�a�͝͙w�ρFXe���Fr���,���Ƅ}���H2�������T�|
5S	Ӈ6���؊?Qnj���6T�^eƝ98�3�MG뙀jI|z:����T��u^>�?g�Ȋ1�ʄ�`\(���C>��#y��y����&M����4�ݕ	��=T�R�P�y�oԶHZ�}*���wR� ����1Ϙ*{��p��0��`l��fլ��l�]��uI=��������z��g��f%�y}�21�p���,�&��">e�����X�18Ӡ�d{JX~͛�!5
��$)CO9�9��|8�H|�M2���9�%1�3~Fq����f�+��Dcm����$p��C(Y�v�q�>�5a��By��k�H���Y�:-
t��݇��V�e�X�48�@�/����WGS��^���S��đ�pnO�#��,F���N�+��l �ʁ�z;��$Oͧx��ѝ�FQ���eH2_YnT�H}���r�bj�I�ڼ5��9��?~ ��� ��˸�V�c}���"T���pt|Ig�n��r��x3!���)U������QZ1U�v6S�d!��&����N;y0a����Ξ~��#(��9��p�pX�Z���؈K�-�����x����J{z��\���ҙl�BI�ݑ/q����e1�tU,�N&�J��ؽ���8�+��40?k��i\�~�YĒ	+���'���;�GkYJ�,�oe�[{nͫ���W��j��"�	����p3�3�hg�Lc�a*�A|�S�'`=�PRJh]����p֟�j���5������FtN!��O*U�iݠ́��F ����٘���t�"�f��u�v�S���**�//�I#�t�sޒ�3�9'��L��@s��Ma���%E>�0L�=Ô�q.&��9�`NT��a��p�z2� +���W��ō�=%9�ޏ9�yR�+k��hi�����;�.�<]K���]S>>1a- ���>�ɥE��M��ն��������|������V�����@���PR�i�k�~7~�!D��"��p|�� )(+'v!�b׹�z��P��0��7IQ���E��aO���T�QC�R2|�0M,]4�H�iӍ\I��[��C���U5��{4]��O��L���Ej�oxve��CPd�٘��:���B�[��8,����w!8#jB�B�;�rD�2 k}U��i�@��쮸��rՓpCp��PK�$���
����!&n/��[Ȑ#)tY֮��1�_W�P�d�K)�Dv�JК��w�mT�$R���v�|�K�,@4��_+�dԗ��j��/�__͑��X^���L���q<_�����$������#�DK�9�!���\�����%Q
&z�aY��dp����?<r��5��I"��/e�ߎ*�_x���)��)�x���ڻ�@�QC�2�����~��4-C$�qө��v`�=��c�=�|(��B����;��&�`bu���E�cS���G3�e�.��8��q�.[�=��L��,h�膁��_��Nߕ�;c���VrکT�(H����Ƴ��V�
�=��4c�m?��gҢd�T{��g��$>#>���]�&�F�D`�S�ڞ�o�p=�ک�\H���5�i|6Y�_�&%\1l���vK�	]��%2�S�Z�F�>�Rx1�䪨<�.�� ��?�3�`��x2�(���>��ė ��d��f.������ȹHJJ�!�|�h��b(}4�/D�L�/¦f�������f*h�y�$����I�=�A�Sok_���'�|��1�����G���)I��=-`��U��+��3��)7v�ȇ�W:e��Є����)2��K�v��b]���4{o;�k�Ε@pIY�]5Sr��*9�3�'�� hߪ�%A����cpL�U"QM(��~�rS.%��ڧz���#��SH���6QD�#=��Z
����>3bd�>�GP�1��c�Q��=Qpj�#���u�3�X?jE���^3�V2��ˡ;���l%�����:{T�h;?$ͻȢޗ���%&����i��`��K�E䴬a!�X$OH��e���LZ�Գ_�\��*fm"޵��R�LLlGLF8o3��v��	]��7��u+�h�>�l��դ蓌 1�>�)�;�U-���.ʛ���S� ��ս��DWCaj���=�%��G�~ D\͌�wUh4rBv��6�{�~��f���� 
�З�V�7T�w���s`��U"?x��m[:5���p�k���s�}q<��/��_�]���x~��f��N���)������%�1)7Nl D�z����<�ļsn�n|�����L8hZ4~|�)LTQ�V__�� �lS��&E&C�=���'+zF�t%H����1�<&c���M"�ho��z�ϑ��?Q�1��"c�Y�N�d����
�~P��O��*�f=(�����_=�@��ݵB*-7�p�Z��B蟎��g̲HhE�|v%��>�N�$����.�Q���u�`�r5|
lmP0��l�&��W�K��
�@��|�����7��#?�o���AB aN~��(��cs-:�_�7`�� ��i�GS��d�t\b�q��q����\$�VƗo샯��fzk5��"��-�����J���4�,&�F�3��W ! �U[M_�\{?%���c�F;�Y7�M&���̎�D��!F=�]��@;��ˀnC�d��l��(�u���7}����;��\�����O>�r��f��KԣG��H�2���;���7V�Ao�1��g��`���MW������_c�\x)��F���{q�T�/?��9a]�_�������)Ô�j`Mx���,*F��1"�Ь�i�4�E�� <��$�	��b���`�2�E֧>�kQ�7[)��Vh@}�
y����~��|]'�$é���	��o���v8�����E_���\I�j�]1�k@oM������X86 ǵ|�O�ȅ�w>L!�V�9̗���N,�
!���@Q�4��X*<�9��(t���j�{j F��㼥�"F��$s,Ǔ�ۂ���t��d�{��/��2C3����?��s����m�v{o�ep�Ҙ0�	VR>��3~m��gP9����Uc<Sw��6^�t����L����)o�z>�ȼE�#LN������@�9�,=�k)�0��K�/�B��Ύ:b,c��CH����a�h�u*�T��� ��{�=OQ�<��nJՊH��b �j̞9�,sp$\�.��*��w�2��i�M�o�0Jf��K�E��F��: 0�mD���
8� �������`x�Wa2�c!Wȭ�L��2GϏ�csfZ^�+����E�d��C�]��f��&�_*�#�