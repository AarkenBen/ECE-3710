XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_[�w�\n�K}:���x�o5.��_w�C��gڢ�;�Ԡ):�fU3IG/���ǹT͈)���˾q�лv��r�B~K
�vP)@�Ro���h�.��Wy�S�*R�zv������fI[�w�/�8��Cn $�?d�E�AD�!`D�-�H%n5�PJ�
�J�R��堫�lGFj&~�?$��zU�ϵsA�!6K�طL�/S_O��J|w�xQM��Į��r��KT�5;�>J�T_h���1����xy����%;-��j��qpN�7�u������^r�u�9L�E9���m�_����?�tͬ�3��5��.��qpp�k�[�< ��r�3u�+X�"$��5�x1*�ӱ�F���ncU�İv��
9��2�E2��Q�������ŧ2���*���B ���E���u��2�6�j����6�H P���1J����ú�֘/�	3z�6la��=��nK9���@xo� 	�L6��S��Er{��"�|�F#��V
�u�\FZF���Ȥ֋��.k9�F�O�0�����`��y�m����v�� Ay �^��Y+�Z�J7�s�~�����E3  �U�r�u��>y�+�Ȯ�8EJ�9��`�7$���5ǔ�NI�׍��Q_.�`0Z�Dq�{�>����J�@�j��R������w\��(t;	w){�z���#6a��蕚�U|0�ڥ��7U���g�����ci�v�QrI�B 6�����;!�XlxVHYEB    fa00    2910'R�{�a�9N-w�9�Y�׺�J&����!�N�H�`��$���'��ֹ����&��>�S�v+�?~�����qR �49�qI'89����+��W�+��԰��d��#vE��7O�Vv荭D�|#%�H�5�ӫ��ɐ�F�w�{��"��M땖|ЦxL���"T������L(bACW��zw��4�F�LR�	���$�>"Wlܔo]j�l�X�����v�^�Q��4�$:�2툲b�b�^ VǷW��q��M��X�,�}�ŸJ�c\��d�]��7��Q�e���I�m�h�R�"dƐ�,v+�����ҧw�����Č��/��]hռ%�BWA���l�V+���t&�
N&o9r��ZKԊ���MeR3����[�*h�<s�}�j����+1=Ι�T�lt�i��s�^d}Z-��
A�w,��j5��Y�L��3��ȀM�'}A�����e�PP�_���?��e��'�h8����(���F�yG�*r斔��H"z���	2�� g�{6��0�߭�!j>~�kD������VEM~#h�]&�S���O��
��5�7���҉`��ֶ܎���12_3���_[l����}(���-NIHJoWl̩{Z�����[X�"�F�.��慆��C��7� v��d#����ɞX\��H�"�x�� L5�	
�(�(�"D�S��GUd�f���f��!�nm�)��!d���	�0�us��ڎM��O���C�K4�dyq��猤(�vfWv.�5G������"+���`P�zW�@Q:#�D;0����I0��� ��T���q.��,p(�!�gF�"�+rmF��\�w��kA�T��d[O���N��.{��K�Ò���vU����p<:�_z��0�W���0�����]\
��ˮk��=i��'��e�5-��[�_me:�� �H�����V*|�lG�?�j�A�~;I�w.�Ĳ�P,9��~В��!$��K������	6�t�f+�>���fs�eM��<�!o�>z*�\`�����������^s9���x�ȟ����魁����l1���O�� ��σU[���G$����-ي\ǡv`7J���'e`gUs�G�Y�R|i2����cd����-��f��!x[% �=�˿y�^I����������R�{(�>� !YՒD����� XO�N�m:�r�=F i��2��4�5q)V��6�.���L����������h�݂V���E�sz�w�ʃ�=� �5����x�I̏���y|��7�z�RP�X
� E=��Y���y��o�y~<v���7�rG�ն{~�+�1dKB�H��l���;o=VR�7��k��Te6��f�z��Dc�X7l³�#��f��+���R��&M�F�+wxݫ��W�6$��m�W�>ƀ�!X3�+��:����$�<7���dVQ��.�����%<,c�:��*�y��SŸ&](���x�Y[�Z�#W[��C.�=�,�{-/��gK	<�ZiB���	���$7ɥx�s^����V��}L�*aCM]��G�J�`�^�"�
W�B�+�� ���j��5��`S��3k*���6d���f���+���絅����"�9��ʭ0Q8ڑ���ZB�l��h;<��1\���buU�m������Շ�.�|O* )4i�-�8ii�����*<��W���UxP����]���`f�e%���`�4����������IJ�>�U��!�ˡ�(t��7ش����?�Z�S"�V���we��E|63O�8:��yO�r78`���&O_͗�:6����]�A�������[���|t���V)9�V�c��m �@�nR3c�[*����12��	���o�%m�[� z�b[� �1Z��2��ǦD� >	���9Li��	F�o�݆y���T�iU2���g㬺��X�[Ŗ@\z95h��Eq�k�
��',Y���?�*I�~���ŗ/ 	�3�^����K{�Kk.�D���L9z��2v��M>���7��&���?|�F)Mxu3�l4�=�ۋ	�����f��5��#�E���Q(�<��Z�y��@J�X�^MM�{���3�K`��IW]���j	��˄{xNfm$�����&
A�s`������)�6/A�/�.������1����̾�,]�?�]�B��dcR���*
��Ù��`�K9!�,��[�64�۵qC�&R���@��XR���T�u]��N>wy&�Lw�n��Ųf���*�,Nn��]�C�mLS��Xy��a��0�qR�}O	 ||���^CK�������u�H���Y�@���z_қkJ���'��PUN��,�N ��*~��b���z��;�g+z��� ���H
�bZ#I	&�$�;Rdw,o))�]�)�V��G���*��$۠6�D��8���1��(mu|=�ܖ4UIk�*�c�	R�j:�����e��R������R������8w��6!�����d��8.2�l�8�֚(JKvk/�VV�JC4�����5p�5 ��9;��pP�����}M�[�^NE��f�N�Q�� �(���y�K�Pk�ɟ�6��� ��"�r&��C+�������� V0�[��Z�
���F�f٪E\�ۮ���
[��dݶ�ZY�L.��F(�w�5o+R+n��Cng
���z�QIq���		��!&)�5퐕���C�G*�71����Iָ�0�7wY"f-�%:�tr�@�F��yc�J0N'��$�Ú��\V��%�	�C����u�d6��"�t�р ҰԟB�3�}f�5k��Ho<��4��p�aoH+i�赖�"���2#����g�5����F�M�/��������q�j��E=���/"�{������ ���m%��Ѯ�u�T*	EY�93ݫ�v�Ț��X+X`����������<� �?_)gj����xr���h�|3Q�N_1Be��ј���/*����s�h��̀�4�������]��AX���O�&�P)�����Pqy�~��ƅI=��	e1���~$�?)���*.�FG�Tu��N��m���Q�.�n
M^�Ը��x2���d�G"�1`sx���u �|�:nh��E	�/8?ɇ�k�_��F�H����K	�s,�
D�͘%�[�|��s�8�R���(&��l�K���4���U����~L����`�U�K��]EFe'M�d���b�3�Ka�L��l�0.R-4����]@�HY�5�E��������)�I���#t�<c�����̐���q�ȳƮ���2��JT��)�(�Ar#���[�7� eUy5w~���>U4��M9����KcY�a�t����;S�w1D1�H���]E�. g��GG�E����ȣ4�{k�4	���"%]�;m5���;����41?}�T�`����+�C��̿���������
��7�b�����(}ϖ)�Ἴ�������{ L�&\����_74� �d�"G%�x��P�r|��5%���ⱺ�M�ތ�"jĠ09U2�/Ujaj�;6��+i����t0��b�����)I�iK[`u���Ykn��,O&[��e��&
 ���~�0��/�E�RS��pg/PDL�'g}�9JK�{�tj1��@ ������� �l ��_=]0��޴��}|�-��Ӵ�nY,D����\&���EB�
��"��>�iwH�)�ɻ�/����n> ��)�8`���ᗷq�c�%,�h�:���VN_�TE�X+PH
^��C�/�`u��,�Inu�q�xb�f�ZC!��\܂�-��(�[�}'P�C�M��c���0, Z /�������.��{2�~w&����V�\�����W�CG �xX������EQ�Xǧ9��Q8mT������_���~�Ry��2�����]��a�m(#�iv���e�ې�?;lU�ֳA�����D�-���k҅#��_�+�ը2�L���f���yL��t����Y��%q��7��A�z���C>�v�VH�S�����|��~)�������ZMsAĈ7�.�++�0�3�7�v��,V�<�V���/ߪ���)����#��yZj-�*���"�.뾔�� �#�d*W|�g,F���̝=~�z��v�0 �+�	��^�~����J�,��s��H^_��:j�r5ſl��ïY�w	��v��к嵋�U\w>E�덫l�VͮI�L'.�WB����@\�K8�}�#iqX��?��|5��]>i��Y��� N���|��71C>0�{�.���a����LnM'��%"T�]���r��T&�`�p����w����=	��a�|k��X�=0�z�B+�AT����H�����Zx*�*S���+��?�.Q�]=�%�5?��	���E�o��5��D&Ih����a�g�M��#��b���u��!����%Bn5���W�=�n��Ё�cc֨�L84q�''��Gl��7
g����)f������j�,x��2d�X茡aF�gtE��	)Y��h{�7�0+���y���ENu��]N�3�� )!�*]ϴ�����)�r2;�� �C����d���ͩ������Ţ�'��4!E�1���*��0��l|H9f-5�/Y2�1��6�8S��g��'��e�_F��5�[�䝜i����N��$oRL�)��#���� �}�Xl�

�Cf����R��^��n�i#X��tB~"��m��)���RM����Vͳ�qD ��CHG="�)�sn���i�	V}���IHܼ=#����^�!*P���l΢���IA�=�>�����Z���{y<vU�H��I�����2@���7�
�+X���;�����+�1$$��r��Itk볨Ea �jφ�q��P|w��)�cq��0��!�v�@ m����q2ˉl�-�Q�U��<�|��+C>�~��$^�c�1OT�:2�ip�W$S�^y{ ɱ�.Pk����bv�!4۰���b(�x�0�X����?,m�Xx �ٺH��jS�sq�>��[��ҏ�}�XTAs�������O��Q�N�[l���&�jq�U����=����M���C��'0���p����h �T�׀�z��X�8P�֤�}������̅-ui��l���;D�p��N�˚����[Fz�d${i(��������
3���(�:T��-��Uz�xp��B4��tK�ἄ����ɣv�`��@����Eѓ�i@��|�>":��/�4��M�M����K��o��
�	/)0��4E�y�[��g�������a�~1����:������yȄ��{VY�$��^�"���6+g�E��n���b�[�w]/R�9d	�	���!�i��h�j�����p�¼���#}}ye!�����Ie�����CU���Kv	�`���o���<)��ϖl���]�gk��I�e�Z���:�3m↨];��L���Gl�q�¹����`+K�K��D���r+�bؓ�-k�-���2����ʯ��hK��	��{#%�Tp���D�*���7�������h*.�?P�<5��Q�F�\�@a4�K��>�Q�e�U�E�m+�)�"]Y�
�D!�Y���aY�fǏ�a# ��\�e#�J��G�{�=��lѝ���M���S��+��g��.:N�}M��r�}w/�ƀcBk9���)�,��H.z�H�Gl�r�z�:���n��5���O�!���b�b��zv���xM������� �O_���tK����
B�}���:�Q9��c��P.,��Q������V���Uƒ�����ē�Z�eO�X㙡��wX̬��z�,[���X�S������фk-�޸����5���ʷgm8�W��'mx	�'ͦ	�u��ǿҧ�?�����H�����G��s(!��?�m�l��o��5�Z*6^�w	��wj����7�64�8�d0M�/�b[��8-�H �8��W��āY���Ն+�x�?���lo����[ֳp��x�F�J)���d�*N�(ܕ���'���)�&1r��i��9����i<�L��f�z/�2]J�G��x�m��w3w���G�AE���y@�H="��#؍@i��cQ=�� e;�k���ِ݆:������O!T93,�ȷ�e��oPV��9��h��W�cH�Үi��NV| ���"�$̑��̽���e�3
IƮt�����/�yjT����J]f([W�jL𻭧}�����u�5f�E8F:�r`=��Q�@�he��݁z�i�6o�*�m\�>=V�3�`�a2�Xlz��`���_)j��[p�?��F?�Z�&�H�<��x�#q}\H���e�=��Q'�T����b��Q��j����O(�Å�?lz�I����&0�\�S��5�����zl;��^���
1mt]ʽ�i'<��U�}�����P�����A|Z� [��w�N	Wc�V�Ht\|������iÕP~hd�vY$Ϥr'�,�&_��Sm�C��.�'!��9�W=�z�`D�F���".�wE��$�q��R���F��-��Z��� j�5G�GE���:��(�I������H�24�$�Nz)�ԩ�	�%�,��}ڐOk�����sa�c���	��&�6U[q)��$�չ,.��D�>��0����F�ZA݅Oi���Y�e��6_�L_�݆�2T�Ͻ�9=�]�:�Ekg	)IǞG�q@C���k�m���|x�zp{�d��J�9�-��.N�z:j.z�2�D�!	���e2�vH��YdA�Va��9��*~�<aT��2�l7�K1��ė Z�+�p�˜�a���+��������<�[ΩW��0�zؾ�v�3��	?-,�LknSL%H�g�Fjڷ��i��U6H��͚�M�A�Q��'] ���~ü9zF*��ɷ��օp� ��ˤC�g�Z�w���(����Bw����F��u�뗄�|x�$�b;��d}t��2�a��Gԩ�q#�1�����{T܍��Ԙ��!��멪~D�C���v(���	jd�V^~1@���Q;Fؓ��{gؕ�P_�[I�)��K��?[��b���8���W��p?���l��uS `�h�d�N��ό���f���O�n�è<"�a��$^0N�����͊ ��k�`��I����Ҵw���e���g����%��`u�R
%T|���V6�~��~�� g��XQ�S�l�g9����`D�/{H#ri"O9�O<�A� �� �B+e�6���	�H�5����S�u"3�A����U�W V�JȜ��m}��� ����ӎ��f7SY\w߫���&2�>f�3�%Ѥ �U�y�j���E��s�TK�}�B:PJƨ�|��KEFu���lmS��I,��Z����xNO;
�R*��*��\M�
0�S��W��n�}V�-��<JkǴ�T���E%ndp�F<��]&�L6��6.�ǯ����`��0�1��O�O��ԝ���[à,N$m�P��y�9b�@�F���#�4�1�����Db������9}w̩����V���+�-��\/�:�����t�E$*�Ҟ�sex��-��g��u�s��H֏��y�V�h]%׽�~t_.~�΁=��늣ч�n�礥���b
��y�n�]w���ΉV�>�W:����_�f�
��A�-
�����n����E˧��#''�&����%��zR��H(�7�G�E���Fg{�g5$o%j�,��A��Yk�<��T-�#dO�R�'��"�KU(aJaΒ�?�"��Q�=��'mɭEZ��#�gKʞ��ƭr��V�Q�D�y'��8X���)�	��}�SG5�J)�&�8��':�}��3/��	�iN��Rm»҇�(���c�������k>7ٛg)�S��fGR����.�[�cON��� 5��,���suVX~3�S�p˺��c��Mc������e�A�(*����/���W��٧��Ȋ* %d�G8/�p?��¸d.@꿺)���S���̗�l��M�W�,�����S���
t7�*==}(����%+�������iH���.[��V��	Nm-gtl��!�R!��}�����y�#��+�����O!\�p��q��Jɢxi��1b�!d�4�bg�Ӑ��f�9Lև'�B�b��#';9\��30�9z����)y�ʹ��`v����g(#^�g�ٞ�����F%҄�M�ܴrE�&�ls���z���:�Q�����Nl���Y�Mc.��SkG��w�S����"x���A�:�G�S*x)̕�Xev>���k՝�t��Y�.��p����K?՞s6^q6����;lÂ̝ES��'\C][����[��X욪+��F$�+�I����$���U�P&���冠=Ry"�ޏ���G��j�4'�I�>���	D�y-�+��ۤ��΍1<�?
HR�An˓z���v�L�hAϙ*��Ph�X�d�V�<\��@8~v�̙�,�Ddz�[�yHj���>�^˶\b2�l�e��[���0	o�Ec���b����s-8m������0��X�$xy5ڗ�-�?C�Cx��Rҁ[����F}�~*���0��W"��v197mI(so��h��N��7���I1ЍӤb̙!��ӥ\Bk8I�E��6u({�:pl��c�3P^��FǱ��a��kuے):J[�(��_�I�i��.�D�
�ܞ?�m���{�Ỽ�K�Վ�\�w�����iݛ$�����Tk]p���a��S֫�b�p�6�fC�hҾmv.Ϟ����x;�:V5�ꩶ�����ƚ�Q��**		���b�fr�2]PM���j;�{k-hb���*	�n����Ƒ���O��un����@GƺL��.Jp�2�����i�)�'���(u��4"kXV��3�s�4��*�C�q�4�;l�ǂi�5)M*�i�v`��[୼<.�-LXE`c�e4��	���VR���������0t�%�R�蓫4�7�BAؑ��mgli�(��~�'����3s�4�1��e�a#,�\�}8쭘At�����%��^��|;yWv�w]�q>kS��� ���$�ĶDS��M��r�ց�� �8�r��I��]��%�D&� �0��2E1���Gv�y5�� ��v���E�Ɣ)LԨ�����>aZ��;��:L���.99��&�k��Ѷ|��O�S}����+|5�فX��O�+P������]`��$c��������GU�%w��P(!�S'6�7A�)�D�ҹD$-�o�ō#�sV�/z�ګ��e`�U��8��ZNo����:h�
h�4o�,�{�ˢ��K������i^RHgR��5C����$R�T���@��&�2� <��6P ��F�MP�?4�O	r��9m|`ܴ��U9A>hӛ��v)(�6�|[b�"�1Rj�*ZU)	�`f�q��,����=������[/q��*0'�T�9;���sԬ��ɡ[�lΰ��kҎ؏<��ß��mʑ �"���>���W.tq��������/�J��p#�'�;�Tݖh��JrO�<pe�P������%��2I�緾�䖯�_	%m|)
�h����@P��R#ٜ4�}��ˀf0�
2~�npB̊vZ�������^�UU�	�$✧,�5?�9=��s*d@��d�������̇c�����XH�t�䧀���5*�0J�Լ����]���Pz!N����#����u�{1��˷�~��o@@8@\��墄�8�P=����bu3�jȎxg���G���z|��Ò(�v�A\+E�g#\���1�!d4�s�KA֕��@ʑ����������A ��d�]��B*�n��=����^$��w��.aY�2�/��(�E	��HF@oIRŐ+F �7�æ}퐁�ݪߠb�NK�ELG���߲�B�]��ьn6D��Sd߉,^���[lbQ����I����W����Z�2�qcL��UX�'jX�_5���(�$t�/g;���;��e���}
HS��
���0�tYUkF/��^���KJ�ճg���4�RD.?����/�.U�+��L���Ր��+�Hᬏi�����p�la�P��E�8Q�t�T[Gw=(\XlxVHYEB    6184     f80���4.�2wӴN��q��R��b��m����G*/�v.�A9���W�zH.�=D�#�OrQnV{�<O��ֿ�h@�H@�O�c/֫�l�F��ǁ@V�w'�\[[U;fj�,��4Qun"��3���,ݵ�: ̤Q	�N�	)V����t��B!���;���������n�
,���>��
��"?�"����D���tF0~��D�IE�_V��gMKm�����갭�#���Ԅvu�sEj=�yU��fe'�;�ϫP�Fa* @	�M��OݙO�]�9�t3�4u��%�ϡ��"�))���?�z�)%oƷ�����Lۙ[5�
/�Rq��@w�X��#���$��::2�0���'� �wGgH䠫��y���<Z�G��&�L5i/j]t������
�$�"�&bdG�"E�Z�nmf�/��;��Ԛ7���c뾜���	��tu��j���s�Xױ��o��:4���)�,I\���k��'C�B�j��S�Mjj>g�du��0�C����xKE9}Э�(�'��F��V��9q�E�:i!�~�)qV���a��x� ������� u��R���x��w�2��2���07��t�7�4,_�Tم
@ ��I�����h��7+�p��.R0n���+����fM�������2=��]�����L},��5����F�t��y&�,|���]A��#s�0��v�~gM��V�]YU).�}xKPG�B�ڶ������|j6d�N[]n��D6^�n�� u�N9�E�a�@a�����8��{��(U'	�"�>���=5t�fN��f
LLa��;�ŀ���z�}��JK�]�I�T�av���2�q_��;�z�U\���y̞���61sfaR�߳�Y�@/Q��	�A-�'����*ImH�a ��
;S(~���q0�[y����Z뛱��I�zμ:� ��E5s@K�_�t�ef^�>��=�w>�Y������cV*��7��>,�b$���S���a3����2��Xe؈S�a���Z���A􈕯�����@�L������~��+�ѕ�vU���9,��7�]��-Y"UD�׼dўk6Z~'pkeo�'�s��e^�@�t�[��̈�Y��'$͊�X�;�dys����a�P�4U�f����ck7�c0�|]u"h}�.z�>��bN�f�V�_´[��QKd��\t;��eº������s0R��	gƵ�Ok@��>T�n���b��>��6��
�<��<��4Ht���0)��lYx=&�|=iGO)�yV'k<�J"'w~�P+J��G�5#���DWe�*~�U��?7�F��f	Y��(P�ΟMR�B�|,�ސ�̉4��P�7Z�sO��"5���?6�]���)�4��0L�8�+���oER�-�����u�%�/hrx���Ӭ�Da�_-���@D��v�W�`9[SB���V"ڮ�u!;nh*��g�r���K���,W�8߬Q�V�M� ���C�������WYr��?��8\Qsef)��a]�8[�h����"����9��vl"8��������F�L��/=�����'����T3�}`?��]��M �[6�V���͜΋h��Wh��^�YNt�ߑ; �h8��F��%����lj���:�F�h��Ѩr�3�o����m"{%S�DB X�#%"�Ȉ� O�������w�£|�F�ᭁ'�C�:nM�_=�Q7�GǿԽ^��"!_ _��r_��$+N����L���>�!팀�\Qkm�d�o�g�0���
ϰ.�V&G�i���fRd�=�ЁX=��G�u�T�]�����je�����B��|�裷F�#"[7i�<�B��5�T�~�d��]��P��F~^�����o'����`yf���yP�t��x�)�!Js��e�X�:��:@��Tj?�Г�%.��<A��Rc�g��z�X�e�V@���x�/'���u���)�%�τ�j�dt���y@�P��ߗ,yj�+��d<�m2��1K��X�]eT�7z aR �
�9D�N���m��_8��M�m��F��X��8$�W<�n$�G�fǲ&��X���PlWO����gA�+۾�H��y>e(b1}LZo�=�t��d��Inso�ghb75)��Wow��8��Ƀ�: ��f�o��zt���h�I�]��9�[av�j�+���&��H�V��1e 
���uB(�Ӻ�� �-�ߢ�C���Q�����\ب�h(�b�k�a!����	`�nT�Ҥ�N�H.��'��9�l��@v�fd;TC~uk���6~w����֙��<���w$���.�4r�� 6Ψ����ۈ)\�W d('c]�3��m;l���7����-��*��>s&n��p���	�7X�4��M'=-�*�&�K�����?�-V�C0���أ/�z��^�VF�V��!E��<�1�׿zo+��M쮅�i�T��f�;�HGvW��f�i�
�QV�% ]��{�!#�Ψ��/Xi�V�+�N�RpD�u�5ɷ�Hs��*�/��q�8��4�[/PK0��U�:	��_���
_^'^��f��)�0��}����KAe���>�PW�I���Y:�I�JA��!e̔8SY*�a�Om�9�ݦ���cl������~A�m���a3��D��c=�����w��f�cTOYúk^T�ChNM&b��vGC��,�=Ӏ�ɿ(/y��m=)���r�,zF��'§��t�Py��a�hr!W������H�U@�E��ۓ���(A\�����ڳ� HG5��y��
�`��]�EO�kLԁ�9�X�QM*��1i�޲�@�:Q���������+Q0�	[h�A����j#�X)h���
ܤ ɲ��i�y qmO�ߔ3�4��.ᄱ������e��.��;��Hx�rZ�?� �g�� }IO���A/Uy@w�]�)6Ѣx�s�8�QH�m{��[��@����T�D�4���,�������[�$�PɃ8V%`꬈��f~����(��(wC��8b����*���maϷ�*3�,��h=�����(������D@P��9<��w���5S5~�U���3� r_�r����Ik|��?�n*9��ݶeQ�Q���N��'�eL|�o���xH��K�Բ�zH��7���/��@C��v ��0X`IA�G7ҳ�w�Ie�V�
���ζ�KX��t�������Y#�qa��y��g��K�*d�I��co�iy	���ng�6�8�=��?�!���cT�ܻ,����\;Ӄ��_�D���}Tĉ�;;��������}w���(�[�<Lym#��3|��.���&�P�^ �6^�~�s��-lY��q�z�j�!�-ˠv*'&��9F�XT�զ�P�+C���#��$���:a�W�lu)$��Ô�=`�Γ��.x�	/<P��	����S���v�#�п��[���u_�k���g/'i�h���ˑ����W�A��z��2�0����������7Q�So�������xPJ��ϐ�t�+;�����7���{D�M�CQ����#���h2���e�����A%��gw��.�jё��ڜx�=�/^�3��7?��Ʊ	-Z�f(�T b�m�>h�f^�<��_5_��
��>.u�|u�e����ةXU����#Qs��#'�UqX�d���~reg�7,��61�iM��A�Ź�e!���?O���F�VFK��]�s��_������f�B�2Mɯ����4 <������E�3�f��s98���#�I���3���NL���+���'�[޴ �kl�n��c��ds�"��e7��b�N���ab�Q��~�A��
��5�E_��:��\�a�������