XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�I\
�~���$�96a�}y��)��D��N�0>=�8Wt�;�>i��r;�ȥ)eh1�I
��>YC]B�uvRH2�������9�c�]���~K��`�a�3P��F��na���� �"��C'0�P[�H��jm���_��:Ƭ�g�pNḒoZ����$.v]�}��gWC��'���¤��ǂh��1�sd�iͣS��d��ĳgNe�������]k��&�i����Wr〵4;�6P��~Z����.����(�۬l�-Ag	cj�x��0�+�x��E�����Y�c���LX\*y����ݾoa�����Lt\�2GN�4�.�]�0a�(x�q2Ҵ��j*��2X�S�x�`�x��g�na/��%��p��"���6���d�b�s�����&	����}f${�-�
���yQ��8��|\���� �p����:|k�R��r�~8d�*{�jf�٠�QQų�j�������bP �	eT:�2��VANh�"�|��F%��3��g��|.�ĺ�&����@��{Q�ъ9)�c�/�.�#�ϥ�%�@���]��+��Rί�-?�.d|�빴72�L�'���z8��5�������x�I��:!߄9�N��M���f���G��ٵ�)��E{�wRs��UɛDoT���\�7t'��	C}^�����el�/m
�dp��, ����G���k�&�I�E���q�۝|t?n���L�׵�M/Q�Y�F5Y�aVۖ&�6XlxVHYEB    3504     cb0?~$��S{���T���w�w��Q�Z�QW�!�k����IPT��
��(j�m 1���1m�oc�tv����X�ZݳE3�B$!iP{���7"��ס��9�Z7v�+>R<�֧ۯO\�z�c^OA�3�ب�B�"�0P^�%wJ�&��P�i>�
W�b��哛\�S�U�u3^�-�uGy	�T����L
�A!��3�0��=%6�?@Fr�bpP���-�E��lZ��r/���n�����_Շ'�Mw��j1^o��X�m(��ˣ��}����<(��F��=���й�y֙3�[��Y�i�{�u�����<�_A��^�	�~��H�-�*��ee��|V)�����nw��-���a�..�?���<1!v�̻��s�Tc �ᕮ��ȑx�P�BM<fiT�*�h8F`N8�>.b轾�������CHpV����ˉJ� 3�I:���<;���z��tqbE%�O7K'kJ`�3,�b�j���\l�~h��Œ�nE�]�qauS"�+��_�xA�b>y۹xM�5�f��0F�]��s�k:y��oLK9](���䌡�,H���Nt��k�e��5��`���s�	{T9(���Ʈ��DjѼJo����ys
p���ґ�هf�-�g�_�>9��� ч�h�*e�[~yG�u�Sh��4	�[�#��k�6���� F��z�h�KT1�<�F+��a��J�HOY�8L������y�,w�`���ƥ�Mv��%IB��}����J�e���\��~B]z���1��U)�'�Δ�n��a��xq�7��&�Q�Φ1>�dU������K�Mc�ayX띪��FL�)Iͱ�O� �ol,_Ƿ�:�`��?�w�����&��S�䡶B���s�۳�Lp��!i������
����f"��QZ���a�:�˿m`B);��Fl�l}\�qW��2���i��?r@2�fƼTG	S4�l�b� 	��<<���0,PhJLN������!�c�,�O�VN�������J4�-T����GQ:;-8q��� ��6b];��]��E�[9��B~in�߄I��L�1K�]���rӋ��<��0���7�;�|����CV���4�C�C�M�|����~=��H.7
�7s�?\���8������7�)��І%o��t��?g�a3m���b�b�w���S#27;���-�y�Zꨦ9�3�r]��0�r��ʝ�a�>l���Lp)5�=y`]u����X�Z�S`�p@,H��>�"G�O��V<���~���4�YH��ȓǗ�~���� �LI�N�wILTD�Lf�+`wsH�a���um�G�&�� '��:�\�­(�w�i|����d䜏�WL		��}Z�k ��EqYU�;LϾ�b��7t�%=|���%���#����\	�Z���U�E"��� ������ ���S/lz�p��~ z���2�BbE��l�}]KiN'/�e(�oe)Àb�s��W�B�N�x��۴d���&;��3D��\��#���9�M�/|}��_U> �)	Rzr��{B�}�}UO�.�W� �D9��:�-�(��z��cu.Eɶ
�����mR�!��֘&��wE2� �z4�V��q���'���R�l�f�I
+�NP�ȹ�7�����\)�[�i#����,���s쉨�֟$�ᅄ������m��P/pD麍��S}6l�n`b�$<���H����.ԫ3�.�xO�l`l�
O��
=&ѽ(g.Z'��ɔp%5�:$��;��;�Z�mT��Е�6b�<�.��k��eo����Ͷۏ2��o�e������.�x{aX�'�%�O�t簡�D%�V��ɪ#�����h�~��K^�	8i�G`���Oe�QZ����lz7�?CN�י��Y�߽���!�E����}�d��Ϭ�
��"��!�"JI���g���U�?�H�	O�?s��WȚU;l�L�`.��2!��,Bŵ��Џ�N;;��&@�Sא�^�WS^{���B�(@2�in֕�2���\�k֡��,+�%���Si6�V���*�X�Z�4��X�æ��zĊ��'��-����+@�b���X�,w��t�x��.!}�+?�Jb��kQ:�z�������g�0Ш�m�>�K���u�t$C{efۋ��	��1�p�y�B��P1��mĠ���?��^�g]����m+��.f�=�g���x��3��w2Nܹ����8�a��QuDE�\L��oD��gy��������C�'9O�	P������+����=7��6�>�b�%�I��:�������H��a��0�$r����.�N��ד\_�1b�L ��>�>�%���Z�G�Ԛ�;v����D��-K�	�FP^�f�D ����"\Kl^�23�Y�]Q2���=O��ܾ���hm���^�9��I�IL�I��]'��SGEbP�V4��2��}��a����xLA���r:%撹��gh�Ƨb���rF��Y��@*R��`g$��%�M��Pޒ�L�y���}���9���qg&���%n�9y��@��4��l3X(�������LF���1����fc4e+�U	�-p/rhl�����g�T=m������&��^� ���Rg�,W�8J9>G��{L��6��^=S�@�{i~uC_M�I�A�7N��bL	��!^�5�D��-��!Z�',�e�6��^���pEU'�̯����R��Wf`P�c�OvSe�q%5Aq`@sC/ـ��+�a���$'���ȍI�ʧ��T�g�߮��#��[�z\x�/s%[N3Hr�
�B��'�����5�4���Ik�I7���TA���C��7w{IOz�+ʦ��8'C '�_�W+�����5�A���c��HM��52wG؏�d�[O�`�s�zc�Z��b�r��}�s8ǹ��8�'(�����m$�Z��3��ߊ�
�p�[4����K����C��sL%KS��r?a��	!w>"�t�6���V�i�.?�>GY�E��o� ��|�6��R��r�1��&�]�G^C�oQ�EoӁ�����jd�bЩ% ��r]���"X�w�I��D�㴆W�(܍.@d0 �k���r��:��eܤ�n�ǚ��r.�� ���il"��/��W�a��Ϣ�wZC%