XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�L�c7NB�j|�@
QT���x�jť��m�Z�7���Sݒ�Vb�y����hT�~��_� m���:��¤B/� �`��ݜ#D�z:r�e�SR��a ��cl\[}�=���޾%y�[����T�k�X:��/RZG^�z�Z}��{B\w���������q����	5�r��$�w!�]U�І-N�T��L��z�����Gi�E��2�ğ�7`�(C�qd�����aI�Jx]�N$Sm�T�~���Q[��E���I	�[�=AR��Ĕ6�����ʾ�}���Y�i	ݱ���儰��Bv���
S۬}��K�89�
v�q�#���-\O�m
�|�%C��Iv"eD�>I�K \���<������WP�f=�k��>��=9�j�]1W�\��~��,�3FЍ?��?�k/�|-G�����QXn��
��֮Ȣ�'��֧��2h�+WDe�V�"��x �W��<>
�5�i�\�O��/���#<X�<��ך�1��
ϔ<�MJ���̑�;��SѾS�b٬�ѱ�7��R6���K)A<�o.<BV�FY�ՙư*�6ź�1腖�W��`qfa�]P��_��!uШ���If�D���t:.�mו�1P��Y�v�k8�U�Y�Fy�*��{���[����Ӛ+s�A�n �*ƌ� d��@����dT��89ӹܝK��;�j�K�f�[cN�T���S�����{Z�7�)��$�܂J��\b�[ r�(�/�XlxVHYEB    fa00    1f80�u<3��ye&�ĚŮKV����Dj�\���P}�'�Y�΂i��su��L�*��*$�Ffl�d�Ҝ��$6!�:*O����
�`�)
�>o����qn�?}J'��0J��mV�JTD����a bh؎����0.8>�%���X��/դZ�:�Z�h\�Gh��� Y��8�	��)����ܼ�����l����J
Ug�gG%SJRe;��z��E��� �VY�K.a��~
w]�8AY��/��3>��U��	e�ѿ~�IF-��u�i�B-u��=���ǧ_m�N��x\!�e��Vލ�KF�V�����OF�c^���sʈ8�O��cޙa�fg�!#g��}1� �w�F��_e��?���&{C,F�]��JO��cCW8&�j(��-���F��AW��MSPt�߹����|���6��E��|���l�Vto�o�C��#����D��L"�����g���[+X���!��8ْ]?b��a-;uYpf�O����f�Й�5ۄ���-��I
%QM!�Wӆ���#���c)�k7��<
7uO�v�w�*]�ӱ��6�2�m�dw$!���{�aa}���ex�O=:��12��\.���q�sK˾�W.o�ޮ��qO��V<T�E�w�Ϥ�=�rVk���@R�3�AJJ��C5��}�S���=_i��V�xX�J�z"��쐾!$9V���XW�'|#���ōpu<��8O1#(�<�8n]K�ٌ��2�P�Y0-0���,��<���%u�Z���?�
yh��?�E���u�����y-�*���:��	m���0�K�-;
C�s6�Ip�����ysi�N�P��J ۉ1A���M�i�%n�#���,Ҫd��9U��Waw"k�~��p��i�� t���`�wܹX.�rW����S���-K�@��H���"���t-8=8击7�V�>� �,�>�����G����g󭞀ӗe"{�H���]�[fb����ר��b]�X§SGgQ)�~R{D�k��j�M�2�k�'),�m+�C!mY�(*��ǂg�w�>o6���`���2$i�d =Yr�M��.6�؈��Ew�%�"�N���^}vt��EcQ���1ŷ�i������H��YB/د_73Uz��!���G%'�Z*����bKtSC����h�ȶK���p�el5�,���܈���[�,i���"m�=L�����Ҋ؝o[��+˵&�W^	Bǂ�G(}U�0$˫,�h�"lc�u��6���3[{�Ld�ɤN�P�J�n���X~���P��ҧ���k�]�
����}
����ww��?a!��ʂ1pX�,���Ě^Ios��wDy�du���^X&#�W�"w�o�:�A`P�Wď*D�Fؾ}?f$�Ǯ�Y���T�>e���\Pc�_��� n�`v�C'@�h+��g�-�f�
����~[&���뺖��ػV���8�:��2	�V%tl�LZ�A�XP��Fe��Ţ�s&BX)�c�S:ry4�@�qf������Q��o@���%��A��Khc���q��>��nLL��G�mw���+�+'�M�&�b�.x�i �!f���̓�]%�AF��������~����"|t�ksw���	�뉽�I��L,j/�3>:�j��o�dV
*#�	PZ�L��b��X����T�t�K^gP �1d���հ��1z�g�'k#o�Bh|���E�3g�b5ݑ7u3�",+0_wX�k��ڌ}O�L[������~ޠՀ��D�������K��,еٴ�L��n)�Nf7-�oZ���جϋe_@mȣ[�[�WW3-^^��-6G�~&'�#� �h ��dH���}��� RZ�"��Κ�5\�f J#��N�"�У������v�쮕Ʌf�fX�Uk
}�[*h����¼Ø��Z�@����-�ZdV6g^�/�]p�Y��[���p�6�<?�5��|r������;C��OS��gp�$_�M��_�4�P3�X�0�0QiGW-�I��Ȼf�/�Ո]���;�U'��V�a-��MǇ�A}$�!�v�l�J�����D�ȼ�@�:V[�u�[�>��~e�~�5pEڌD՗Sa��ᄈ	5�8};��+�U��r�+n566'ٔD� ��J�pɉ����b������x�F�,��O�\(z����4h����?:\��T�?Ӑ$=���!ǣL��}Lƙ/s��b�K��;��S�+p�� �Gs!BN^��6)R�B?4j�*�W��S��x����%�H�O�.����3��|jJ�~��M�G�Ieh���� ,7iW����9�4�ш�1W�P�w��@�-h����3�<`�-��[���Y���������c����.����������%��OVX��Hl�, �l>��уv5���̂�"[&�H���.�­��z��ڨ�?x�TG���MI��N�J�%0U�.�����wBb�[��Υ��
�S���� V�lI�4��w<Տ��P"���a�W3����!��M�&�%�E#/�_U�������#5��=�I+�[�� ɞ6$=�Yf�l����[�� T�;�q9�c?X$�� #ua��?�;0J��)�=�z�lRh��vq�u�Ҳp�4T��IGng@l�"�M�����+�n/Ct��7CO�n���z��+|x8�������2K�% �5uȐ�5��賩_/3�ȼ`F���Ű-�)�C�=�<���z����J�.N~zQ���3�zw�0Ь����^�,98�]��܈\��p�B �x��Ѩ�G�=��C�IOk��yL���r6 )v���?��\�T�&�n�i���db�@�1,k��E�rI���v3u��GH7$nC�Ue;ՆF�N}kʂ>�M��p"_ޮ�oZx���N`N�< B�	�Me�l�IE�]Z�\����j$1��H��K�� <���4	��Ez�]ҋt�
��t���V~�k�T�^�H��#vVw>�_f��Q����:"�idr�	����z�>� �_�L^CA|JO�X��E;޺a�9NȚV�����p���L�D=��ZJ�}`F
��$�3��i�Q�r���V���m�E,3�J!�|����7��P���	3'("{l$��Y���eCYع���J)67����5yt� ��1u[���n�-���[�a2k�e��_!�)��߅P <��<�'`N��P;fn
g�C��8	Hv�/=)̨:JbB��.gP�����Z�n+��ܤo;[�9/$�kx�N;F|V<,2�3��DA��&Z��c˰�[e���x�1�]bE�;k�8���/���ngi<��̂"�g��Ҭ�\d����6�'�$����Σnf�z)�ќ>���� �BMh/�9X�e͐T��#�o#7޳�ZL=��Zs���������͔���t�ь"v��}�Z,��A>�%[g��=��d۞.�}��l"P����
�~�Y�(�6���I������혈M���|�%��y� ��<�}�Nl*�PW���EH5M�J54�˺<)�z�g͑]�`��[A��Vs� �� ����R8)�I� �Y�(�3��!\G㧿�6���SZtx	��u!c�>��A^��w��k]�^�3υ�Wp��~\��b#]�(@��a��w�95�0�,��]�d|��x�IYP�w�(�(�ڌ�I�svn�=���싩�� �9v��U�>��O�56��'Ä/�+��p�"��z}ιhK&�ʵG\XUAmS�Y�""#���3r%�	iptH!G�I7��;O�Y>�EW�1�k���`�`Wb0���̹�H�ݒLm�;�h�x�ܠy�3��P���f|��PL�ͽ���.�jZ3�v��R/*\w�Ns�����`�XE��Iyl6rF�7��*,Ҕ5�U��(���� ︛�v��%K(G��x����,�c��]�w�?�����:q���=E'�ߴ�P 9�x����0z`)&vq��R�ɹ{��e�G����N��� ����/��$��/�M3���#l��?��݇BjO�~`���1O�g�H�F���a���^jNM��E�#/��&�Q�Gd�?����0�SGB�Ft����?�M�DX�|�� l�/��p9{4�8��{��gA�bD��}���6]��Ӧw8#�V���nC���A�V3�C�	��,�E���I�*�>+�[�̖�(��)�ġ�UC^�3G{M�	�Tu �@�Rd�օs����¿�T���2���-Oenv�����6~��H�|潍QO��>(z`�?�N�Rۦ�+\�K�^�&����k>�s�f���gnn{Ld���4���{�{�������z<�z�z�����ұ�2����ʝ+^�Q�7C�~W`�J'1%�cJO�����Ȋ���:Y8צ5G��IK3cE
���%#��N޴�-��nfF�,�_y��x@j̤����d��d���6o�r'��x�[I��lo��~�����"��Q��%���z�S��r�qID�B�Q��|�,�j���.c�+I䦺�6�R-�uX�1��J�����r�t� ��������4��d\Q3 ���h�#S/{����4U�vc���\ꐒ���b)m����UC+_ T$�/�c ��/�g�)�0��8��Ե��y��~j���d�{��ZN�[�9��X �, !ے4����˺�T��"���WEf ڰ�S:��D���5\�י��Y���޺u%���>A�w� ��;�^Z��؍���*�3&��:3�R�PۆZ�cB��l�e�%�&���c�,���Rn�/ɤL�pE�[Ĝ��L/M�&$�d�=��L٤g��6���~ܸ����O����l1D����Aݲ:�O"ZYX�|���k鏷{fîN/J[��T�(�{�5��Tn/�XMs��ˆ@Z������g���̂,�I���r>U#���C$~>��y�C���Λfi�:�l�_@��i��X���߼�/�fE�����Aj�$�E����?xL��MW0�cN�&Q0��0�&�!o%� P��l����B!=����Fm�-D�Zf9r	��*r�=?=1kW/��?-�0/���Q�عn�ji��SBі��{�P��c�b#��*�)�z7�cp�6tT�����U��$�sA��H`�_c֘Uȁ�1����S'�Vd�h-�V�r0F��(�_�$тw��=���<`?(�6�3^��q��h�� �b#J>o��~owI�BןJĹ�? �t�1���o��Jj�Ol���1���8��C��p����	 �Y���Wj�aU���b]�lK�Dw��kp�0�����в�=_�˞����i��c�3(7ca�RC�̄�B����|>q��F�E$-V��{4Y�?�O����xJ�Ҥ
���u�p�;�+�@��5�~8�\p$�D'��Bln}��Z��W�����8l��E�B��~��CL�t�E�U�|=��ext/M.
T�o�?�$}�����ee��x&!�0�h@��篑+������LM�E���r%���I��q�����o
��%0X-xY�E�i���;�����BR��������?��H�6�W�&�+�h��8��BA3�V8��!Ӗ��0����;��w�1��D{@�I=댎��p#�V��W���l^�'��e [Be:����Ӄ{�}�&��f�|�jY���$=�g�	��J���*�=��a^SY�h��h�M��og�٨8�QPi��P�v�?ғwV��AМ�����+5e	wP�݌����;{V���@�>�N��W��7坎���v����OZE�&����9�0P�%�_�tc�ޓ6c#�+s�δ|���%�Qb�\��š=D�@�Y1�-�j*�ą��R!�~�3C��
&ěL��ü<Tgn�w���8	[G����# Xm����`�hM�V",R5&D�H���L%j�1�b�˪~���1d8� /��w`y`��x�v��Kv��6�o�~3��aa��D����J�(˖4�'����yi�N'�B��݃(z��E�e��v�@���~�Q��*��Nl%��-2�ǵ��i+�����
�Ӥcӎw�\d�g�ܻj#�� w��X��XM;=kG�M��8�wy��>��A�)F�-۱~,��zk��x�4l�>�
�L�v���S�W�+�"0B���������B2�'\���?�M$��N��@���t�x_��e�ں���o\z�P�	*�N�|�����8k-�D{V؏��yy(B�Jm�r��&R�.���' �5�#�!��;5�Qc�4.��Lc�����գȎn��X£����nh�Yآn��
A�RC6H���%��$�F�dJl����J�p��
�\�J��n��P�4b��d�4ȗbM�t�� f����bڊ���̞`"����H�Rvh��W$ӌ���ej����z��"��~|���H�.�FȠ�����%�8G쭼���'09x�S4t��kSxPi�X9�!������H����:zX����t�P�I�-"�F�c���U[����<�Z����C/�=;�R���o�{� �<��)���������ӓ)qnF}�ڷ�p0�y5�"ſ;���%q&������/K�=Fi�.�<��e�tr�y�����E�ދI.�/׭,łF��ަн�	BN6�p}�� AQ.6��𣝨�w6>�����jXN��^���ȳ�U��Px��M N��9��[�q͔�M���M��0�p���'�n����]Ct;��S��>hg"z&�<"S�kL�;J�"Y�}zפ2Z��A�I̸�8u�z"0Je��(pBH���l[UMlrm���H ���\����,�r��W�����ݘ����2��P�:�-`k��VvEs�	�5(�q/��yy���PT,#�������}����J�Nt �UԎC�Y�����ದo�Q{��i�iY�����:�L�'&�$op�«��6�B���1wu�#ߋ��'f�D�V�P��M�V���I�g+o���Z$�=qC_m�݌��#3��|<�>�RG<C��a�t8Ն�s���f��G��|�#��\� �K\���O�"�h�.ꌵш�d����bK�	=���A������}P�)I�g�G��?0��A����J�ۓ.G^�ʛh�$1x����f���J7	��b��UH���(M�#%,vX4T��$?><$dYDD!�iZt5K �Pn��M����d��I.�E���KBT�ۦ������Ɯꎗب�vH����qX0@y���ٙA�j2W�,,~?í��E x$#/ �(N?��}R֪�ӎa��G�7ȍJ�N��t�P�7�p�����M��I��T	��l�1O�؝�>H���Z�io�!`ﶬ���zJ��c'2�dG��V@{E�H�Q<�fv�_r�B���XkeBK�c�)@B�Dxg�)�����y�S�Po��q�u+��&����"ST� ���ISÊV�#���O���M����ӿp@��9cC�|o�zt�������`p���ߺF��gd�(��l��J�q��,��ݱp�˰���qUA�X��N��!|���Fvh��w�n%��S��B	|��w�u/��\�aLC�1�3���g�@��[��˪h(I��C�)(%'������ �{U ��'�9r�e�Rg�.�n=�'j�d�Э���R5��knB�g�V���\���l�jT<�:������!���U,�$E���wQQ��u c�M�q��vvX�"G��(�z�.���A��1ھ`���Rط�Ai��aB���M�o������ /Y�<,�F�94���I���S�NR/��XlxVHYEB    fa00    10c0�-�A�775	y�ZWw;oyh�hp�?}w��##K4C¶f�4�*�*�,6.�	=Y���%�Q�*����r<�X���D;���&Y�!s��.�q�����������f�[�Q����D$�Є� K��腭���L���RH�§7p��͏s��h��i~8�d�	�;��:��W�Z��&X�������,+�@��cCQA���K1�N:[��ȼ}�ϊ��?m(�I/�}���.�b���� �N�7f��9�+0�#�h
VhD�f�P��ڍ�Ơ�,�c�Ę\�`�X�}WH9�)��F'����ǆ������`�x�А���`��6� E&�W����ZѨ훋4
 ˽.5��/F�ߔ��){ �~�pbǉߝ�ӓ(���_�����G�eB�/�#����x����ýD�?���0O�f�6���W�
,7e)�4}���q��c�_\�t_� ���&&�<�^L�=�ny�E�qJ(q�B���.&��x��D�J��u�+�p��Ȏ]��{���e�%��I�Ի�|�YQh����4���9۰1ˡ�W���Ig>��&!Ƿ���J/��2g�/��L�7�R�8/��BƎ;���'�4=a���hVNؙ
/V��q�+��W�/�&ȼOc�lz�\L$0p5�� �s�h��W�wR�t��
mց[ڐu-alKY��Q͢{�87Sa�/����F���2�w9/i��҈������g瘖"�H�^�z�=��ٚJ*��13�cQ��@SV���Ս�Ѭ�.D�s���k�;9��(�� й҂�v�����[]�v{��-��^��	j��])���{;p	����}!.	J �M��+��\x�G��Sj^k4C�0�j��	|�|��p8n����X\���y̟�?�F���FW1w��b���	q�ot���(76Y��9��!�sN�VQ��M��}�!�K��0��cC�����4
����d]�f�u*D耮��I]ӂk���ͥ9ˠ8-�5y#ԓ�J����18E�������X�4�����7|̳_�?��y'F�eѕ��c�cn���#��2&KS�y0����PM.��^����3�#����֐3�����#�"��gx:�<��-`�r�<�Q�n~�M%D����9req��[�\�l���ah�� �ӗ�-�� a������l��Nu��kp1�S�KښoeM��?mk8JH0&��1pvIw��u'��-T���t�OP�u�'����FY?Ӕ�*R�
�:���]�]�F촸|(�Z��l����������l��;���\/�{���ݐ#�9�w�ȷF�EE��j3Ne=�%�d�D��ZE9����̚�E܅�Ղ&�~{Qm�3]��UE�:���4b��0��h�U�ː���^ʔU����q�[���E~х:�����!�M��iP�-��CRi���}(��h�naᵯ�QX��/y�Ns��쟳�Ry�������<\�'r�^�7�$� �.|�m&��ZX3�zG��cvSL�DCT��Z��ߢ�A�w�۝(�=���<�A��I{�2�6����;��W4����l���o#sh��'��DK¼��*�X���_.v��[p�l����A��%/��"AjRx���{Q@73V��6Eʀe҃	'& κl�fY*���/�%@�� ��]����ܧY�c}��J~���+w"�1���j�21��rDo����TZ�p��L����FdU�Z��M�����Rn�{��_Zi?a9�n�T�����j�Cǲ��a>���y	��^W�(vYhڂ��n���~Ӟ���Yy;�=��X���^��V���"�/Q����	���{�d�x�6|��?މ�w�qWo~
��*2(���e<��+W�������]S��{�+@eOj���<7�S����x�<'tF�f�*�r��T�dЙ��E�XSY�͌AwY)�h�ɰLCm?yh�i{�����A٧�Dx���k��r����B'b!ڷ]GL��v��b���~R�&����Y��x�y�;���iai�<�g"旙9���o�,nf�1����<3�&�u�^�����$�GHtw��㶃֠)��¿UNy�����DPR��Vu�!�jhAş�,T�D��ܳ|�5�	�G�'�|iwr���Q�j�z�r� Q�}�'X�c�z���"T$�yuA�I^Ǆ~Ua����rXHѩ��.�8�O�*��T�cJ�<@x<v��v�4�M
�=�����Q̀��"�]~��1!�xX[3���^�'AO��9��8��w��E��=OJX�l�ql��%0t}�\Sh��C d���d�g��WQ+_��J��I�i
A��e�kx����_f&�d�5ф/q�Ke��t��%f]��C�4V֖��*��be΢�\K�<��g2X7���&�[��H�^wS�A(��$K�|�SA�i���ޤ��=�+6��q��b/70�@�xZԸp��Cg�.�8+D���jU����U�Ek2�,�-5N���d���ܨ����N�x������������c'ܶ=�QJ�?ġ��'ޱ9V�9s,qI���2F�8���裚jg�'*N��܄��o�3�&�ΙQ���^��9+�2���l=�ʎOR%�%D1|V���=��)�c��e��xy�ţ�A��\G-�x�-�f�b����6�p�Wq���mw��zs֬�5�O�P氵N9��[�ᑚ�*�Z������^f_����}sЮ]��W�����+��;����c���0NC$�"��l��X�}���ئ~o:���\�G�d$�W���,<TV�[s1�с�:���(�s42���#Zy��o8!D��˺!�J A���_�3>�`�\IS�+�BWI�R�V����g�I�J��oʵ�œ��B������E7a�#�ڋ"wl��S���,xZ4��1��<�Y���.ɲ<Lx��sk�/=���P�y�'���qX���ɮ|�V2l��t���g<�x��U�9c*�������1?N4o-�6A"I����C���~+K+1�o�m�Z�C;�x������ܽ�u�8�1��XBQ����"x+�Y*E#�m�M˷%�[Mj�7�Cw�c ��o ��7<�t��><����W���� �u�e�fypq�6��y���_�9e�G�&���(;�����9��д��ĕ\c�GZ7�����|&4H�P�6�����*&���%���7��o[��NY�yuD�8B?"��_!����2�jD
�%`�h�`�-3��rz����-^�HI�|��N<��	����9l��o�W����/���cXSA��y:o9�Y+�>m�ܜ�a�5v����%�Y]+RI�o�-�:��?J��h�Aɡ���A�5\��U�wo5�����n�Ħn`�ƍx�˥\��bs	 �̚l�o�񜎚%p-�A_�v��������)�a�j/�����j��\]�v�\������"֟�M/�-|wn��,�M�v!�[/��˾R���°M2DM}��*>e9������ݖ!�P;�W��d:uо"��:���D*�����^������>��y�_��@_�������/�f0d0ŋHG�(H�GjΌ#���h�<;������^�az��&-f��%�u�ڀC����dQ�w.+�J��a,��9�*�����
�`������R?&X����j��� �Q�M�]��D�S�.x<Djybho4����
5��$$͂o�	j����2RoI���KrAoN�b
�����t�O��g�����f�����t�^ӹ��2�^�����{��<�� �؝MhV�A��Y�3���#�Py>�Sg;:���mBV����6k3Ee=2��Ezk��Y�Y�$���2aFQ{k����|�� o�= �
����)�b�"wB�y.RP�a\n�լB`�_ ��L/��Y�@Ǖ��1Q��T�!�]cYZh=��ub�w�)��[�7ITU���?��,���M�SG~�����!H�fc+"o��7ˀnxr@�ű�iM��.?��k�����p�v�fc�4Z��}�;v�O� QL>�r��32n5E�_}��_|���"�NQ�<zq󿎻�Eq��z���ʨ�=��,�g������Q?�_~��I�ą�W��1<��ޣBy��#�?��pǆ��d�`IQP�b�̘=��ȁ��Ǒ	��*v���k�XlxVHYEB    fa00    1140����^��֛hƃ�]��?���U�i@�[���?Y{�Tԛ��i3U�׈^p��=�f;Mb�J�7/@׎'9����"O�ID���j���������"x��M��5��Cm�Zߗ^�M�V�F/��:������4��E����ov/�@u�)� ��9�����	�Z<w�E�˔����!g�PU(��k�=2���'�6E���1G^x�����RP%�,楺��x��J��%矜Hx�<�6���_��	����q�������Bwœ�8��ҟ�C��#M�r�p4AUPNw���@��<��+Y�8���]�T����>l�'���+�2h���5y��lCo2��'O��u^Ci�Y�ݸ�n����/+�C�_k�������`��L�i=:d������ڹ!:Q@g�d��F�6jt#��C�h�2	��LcԿ&��D�/�~y�lp�(b�G����mk�u�F������[S��&���@c]�qY^x���{k�	`-�+o;�µ��<7��i<O�������s��"bs<y���x�3�-N�����,�B�ĕ�t(}��Q'�F��nT �v���<s�I^̔2 �
�Y��d�9"�L�gP��e7�sae�1�D�t�B U��k �-q.��f�d�����oN�vy$�u�v͒�L���_wP�P��cIj)D=�2���8�pLC/Ѫ� 6�aMe,	�6�pƨ�/G�hPTQd�ΐ�3�>�YM[8�Jq���b�M/���9u��s�t=l�B�9��pT����uZ˖�%B���Dm�22�7����(iy�Ϻ�-r8��m��Ĳ��W��*��oB���bc$���ç�_���5Cv�#���?N��!
�P��os��Au��
�(,��ފ9��*:֊G���6������0�˩F<�-��z��m6����8��vy�%<9�O�0��M�SV����Nug�]�
��T;F�k���ߴ���Z�M݈��T�cM�h�ʾy�� �gT�����c s/�:��=���X\�
-D$8�0k�Խ�;&��Dn/,DZs��׳)#Q��	Kҳp�ݟ"��]K`&#�)6@�A��p|K��77g�Y�/8!����V`��*�l��d��\1�$��Z_� X��2���OP��B��D/^�H�x+�Lb�<a�m\�mE�`�JZ�eѬ��P�"WF�g7&��U�]-xq��_n�ͩ%�����d�fW�]��%���)����� ��?݀)#��+�@�[��q��}���������;_E'����$kyF嫿WO�z����L�����w�����'��7�.���X����?l5Lf������Eg/20�v�-��i���,S�qŒ�hf(�k������߇J�E2�[c����F�첥-X�F�<��p�A���g�1�]����۬7���qG�E���9��I�۾�<�,�$'0��q�����������I��4;dvlqi �[���ѵ|�qf�V?���3�*��ј枎8�3"о�צX��]EP2���M�]"1�ȧ$m؛�t_ꂌ{��$��o�W�Ia4�K{�>#�H�Q,޼(AZ������U��	��Ou��of!j��-*�a�k��%�������Y�"Ջl�2��5�Cٳ������[�����Ɍ��Kd�8��������kI*PD!� "<���
�C^O��f��Q)���T�,��%�@��LDz�Qucߣ����{y��Ui&�
�U�}�-��O���4������l� ��S@�\���ҀOˈzD>\
��2�Xs��o����R�8��Q��P��cXx�A$�z�(&Y���+N?ਜ�!aNY�VӘ��w���H��`!��m#�.���c��(J5`&� �B�]AM��]���/�[OW���
H�mkO;�^��k����۠?lW/*? 
<P�U��g��p#���JC9:wz܆�4��j��vt�쥁��u���AOʟ�x�,� �uj?�.�D^*�z$����4D7ml�ߙأ��&�@g��/��f���W}��C�	�2Ԃ�&�>�����j�����R	��1�l$��X�y�P��G�k�!C���!HX�� 좒�Z�u�@����G/�N$TH��XTJ`�&+W��<��h,gE�� _�n��e�����s�񉉭+�������͘	mQ	e�(6��`Xo؏��3�ګZ��d�g�����c�`�aީ4`-��q�6�����6� (@b[�0��=Ro�rI�\;mHؔ�zd��Ӧ���b�2b�Qh�OU*�YC��vP���
A^3��a#0�&�r�%�BO��-�bݽȞ�4n�L2.�����h���2q��)�Kp��S����Me�p�u�7��̔7N��E�]b�RW�(_�]A�@�ZE.T"����x\]�h�q�O�p�������G������E�V�?]�����Le��, ���1�Fͥy{�yC��[�ȄF��F �@��r�1:V��cs��7�^�p����p��3�yxI��! ��g�����o�"D�Fl���#r1�s�Hۿ�Hδ��H�y�U�SF�k�gC�Z�#s����C���u�)�+��ơ?Z�'�� ��ǂ5s%,OL��z�0x+�wu� ��٫ݓW^"d��׍�W�%�.��z�������Љk�z�����u�i�J�f"Fa�m��\��_yǢ`#0ԅ������dI�O�[GfA��yPa[S@x��x�ڃnW|L�i��NGY�
�ɇ\���T��Dq{��G�<{;k�5�Ŷ0Î����a�j��K��6�V�4iK�P~�W��b��5��ςy[j�w�[n�E�i5ӳ\N�@��/��Q�W��I8C+2��!���AV�YR*�äN��L�|-(N���#(�JV�3�2A�JCA�$�I�v5OR��/4�A�	=xK1s��8SxPʳ~���Uj��8���5��G��!�?�E���Q���LA� ��`)T%���4U ���åˤ0w6\٣B*㗸N�"b����/��9ٽcd����,9NoE
�1��%��0.A�pD��}+�j.��IH���lU��Q�fS���Pr�0z�L}�'�Km��E�>�Ge4 hGgFO��!�]��L�E�l$�H4	h�
0���y1?a0Y�L����@�P���<0��9��?��K�'�oc��ӿ�S�Kx�L�[��jq��M�����	ʊsĮ�ڳ�+_����6m��A�7�Z�����ňl��W��Z�U��"�qgnvdvr����gpӿ��j�1�Z��F�������A�Ju<s�F.9����Q?b��^�s>���M"�=G�N�
��م��{�0���~Ѡ�0���1�n����Bi7���6g�Q�JcB+�	#�:��)��(Y�Z��g%�7�r,J��˘�w?�3��8cAE���%����O�Z~�����f��m�V���_�2�?�o]����;/N��F���Oft�ݢ��dtV����kO�&,s�]&j=�>��ƞ�H3�gdz�-���� ���龘a�|��S�,oN��n1��1�J�:��o~z���dA��P�?C�Up�sT:�M�ee�
m��Є@��`�dYU��|e��z���kM`q�c[Qo]YE0ć0�u��lZ�n#�I>Ĭ���f[�C��㿪�#�rvs�'okE<�P�B�hm5v
�#���L9�N%��J®ʡ�C:yR�<Y��m2��H$@��"�M���=�����d �m��x����~�<S�B"�`�d�|�j%5�� ��z����Iܴn�t�*lj���JC� �zT�>��9<� �C�
��yp@���<���Nwʢ���NV�B��C	��� ��Ue���lJ���FTrU-���U��7�1��dP&u�����a��@���6N����yqv�Ǩ�17�+��w�G	��:��d�.q�#1t�B��1L _mzr�~��B>�c����4]��o�kЗ�7g��CXԻ5-l����#-�eա�K-/��M�.���C��:ފ��Ŵ��ߖR,1ux�7����C+.~���&��#N'�X�/�C/�� ]D �H��أ^�=l3m�X���*��g����{C�y��c1���u�����Y�:�]�y���z��v%�Ø��ApLf���$
Q"뭏͕K\l��3gI �_�#�L)}���!��g.���Q�MB����}����ޔ	�`}r��R�2�VF(�� �DK�Q, 8{D�+�T��Z��sK7{]�,F�2:��fV�ù,9��g��Q��D�ͼU�D�/�Z�RXlxVHYEB    fa00    12e0;�c�������b|�*a�jҶ"��F��i��K�l)����z����F��u]y�~3\���	������Q>�ā�@�M�a��K��JmU�t�'C佲*_�V�\��]ː��c����-���(3o�0@���yJU��K��@�Omf ��<�������-�S�q���I%��u�ԟ���0<�0iR�O����� ��%Q�!>�S�<�fj��!�:�A�7"����4��SaUw㧍6~�r ?6mH���MPv>SJ�.�kɧ�(eÛ]��xQ�͚��c(%�I!���%nk�(��E�4�"�l0�4�Hws%E:�����MbK�s�����u�FS��ߓGkY7��������D]�!c����0Ư5ė��أwv"[OĊ(fn#�ۀ[{8�<�XA�����0	���]�cȋJ(�������"r�����`P���V��n]�3|D�r��>%t�LVR���]��H�Q*wK�"W�h5e������E;�hȒ��=��8��|��Jͳ�"31K���Lv���߾��/Bpqn���x�����.�ո�b[��y�፣E���j�'�ӌ��ɋp���J�	�ϛΉ�?>T[��l,�ץq��p{)���VsxQn�^h&�<��qȍ���c(PA��\ ��;��i���t���5q���Sh%�e�I�&��F~�⠂	0k2UWH���+�'iN���%�
�\1�1��N���$�;<Gf�ډ*Ek����3�cKoZ2����s��o|�z�ls�H>��\�gAz�|��+m������ϸ8q$qxJ@�B�qq(�&=�@g�(I���)����"�l��X?EpqO�`a�T�(�����UXؽ���J?�{4`lTSĒڇ��``ߡ"(��#M�*a��Z'8� ����(�(�:G�M�K�&��o

8Êg�D�;�:]>�$�CL+/�f�&r::ҾI�.B8��_�Ӭ��Ll��gXa�<����)������W,S,��_Ya��k!���X_5����e��O	\�,p�C�m�;��s�-c)�&��N������Z�f�i���)]|��G�#�8+�(�,���Y(�d&�v�L7�4��uUF ��j_��%�AF*y��b#�J�NP�+���  �X� jgZL���K(g10������9�˫ӓJ�5D���A{�ʆU�VI�0A�[�_QH���F��x:n_x	��bFI򣢭p1�0+�k�E�3��{J�]x�3q�+m�A� [�W���ey�F��Mkpb���59��A�0�Ϟ_���QÐ���f)3��p�d�g�'%����@r Z�r���?��NqS,��"}�y�k���9� �	�S�^������������G�=��%��>��̊��&����&�U���ŷ���l��6��,��L����T���.�6[�[i�����h��A���b���,�rm�:�w|vv�.Q����[PMtF;�8�{�5�L ��ʅ���{����<C?��$9n����Q���&�dk&��C�2Ze{M�TP�L��ˮh��;���Q������Fv��������@x���g�Ø�ڏ�� 4��C/9�
$+ã�E��5H)������p�?S�o�:UKP�������[!�%�X���c�n���Y$$x��u�Q/ʑ�2�}`�ZсP=������.��C��T�m���px_�O��l[����r[�� %3��g���(�[��j�B�����[)��9���G��9�x1hG��J�����q��&0�
�vd�wTm�a���,��Q��(�Z��@M�a�+��c�q
�օ�\���<#Q=�<Uɴ��u�;U���?�xǎdE�3n��}i��4��qSRY�K7|��g�oy�|���U���ķ<Ƽ�P?i�v�v�� 
��[���*o���$�����]�Wja^Vz�P��b�I�u�D��՛��dؤ�m9sT��<1�=��f����=�J�g,M���5��k�4-�b���/�a�YRN��$ut�����ن�~u��w���E��ս<��l�Ϸ@;}�7Ǭ��zʤQA,�rF�Q����U@�/�&`�W��?�0�
6�ѥ{`v�E�B�`�Et[-L�tE�dQj��ȭڭ��&�Dt����״49ڙ�H��Ϝ/��bA\B5�֠/!�U��o�_�gh�]otP,$��PDiҽ6s�)-.�͏7.�}�B�q-�)���op]���*g��^+٬��	������r�;3v���@Y��1��Wp�k�M��o����"@�f�[K/��-?�U9p���|����	./i�.(͊-�v�Q}�}3�[C�"�yt:�������4���eLuZ��h��@x�)�"�؃������	i��[�8���'s��=��am���;����*��ܱ݊a%�+T�9%�M0L�jH=��ջ�*�Ux���2�lT��T�k#�޺L�ަ� n�/��J�/F,�Ln�4V�Y�IT�"'w�k	�&�SL1Yӝ��Ø�����eN;�(N]��X�O�v%`C`�Ɯ��c�$ �������D�^(�̈|���e�~����ج	���P��4�"���q�4Pi�:�?6�s��b�_oOE����?�0Rmһ��yv�g���aT_{�K�D��u�+�ņ3��߂�iJ�u������L���-R@U��+��V�h��<y�Va
B�<E��!sδS�ʔ�=���Q�>���]�I��)��n������tm����VދZ~�}D[�ev�� �A�ƽ�n�\U�����47�얛���e@���<���$�5�2�ׇ̅4{�\yßZ���/�]v��.B���bFfCa����Y{Zgc����-��?�\��Jդm;V��	Y�q^Rϕ�����"��(�ٸ4���z�D�_!�"��Nw�RbY�l/�ep�)t�����-�YU[�$Y�:������3�qk+i=5P�u#���Z�ǳ>jMt��X7��1�9�����u �mh��t���L1�`�G�$ҟ�\Ų�Ia���
�7?;3�s��nN~���S {n�ר��m�@k[5�c�`���~�ii�l��K����X�^�z�8TE{��}�\����8���a�[U"��Ze<�
���9Q�q�,��n̛�Vxf��pd��D[n��H��?���9�s��Yrj�'G��u��a�;}�i����EKD(s��}�кw5;��;���-� ~`���EdğJ��郹���4�	s{���'-9��FR��6�1b�#�S�D����*��
��h��V�w�oWҸ���rh��4�������Y�������\��M*N�b���o*���g9;���
��Z*}T��n5gN��c�h1^򂾡˴��Ʉ��*d�i3:��	��S�J7_{���q�,����/Q�$ϋ�7����)׾ګ��~����3�����/ *CX� ��wO��)��� y�]t�[�}�3��<������!wI'�2?� _c�a�7e �g⎲&+}��V�����TI{���������[�9�����'4{�Ǐ*��9��n��⥠sU��SD V�Hr�,����C�slS�"PM#dy���2p�!T�3�QC���^�@��s+�_��G�;�>�Ii�z_�<��y��t�EJ>��_�%:H}|B���ڏ�E2���6Ie��+���TK��ةtR�Fٯ�������x��@HW��@��Z���҄kt^��ģX���{�S�wmv��S��Z�B��\�,k�$�m��̣e��?�K4
Qc}��JXa�b/��P~8�>�\��tׁM����\2��x;��d?>�ە}��<�8���3��ml�ќ0 =]I�E��y�?Y���=�dc��aF�G���eB�5R/u��1Mt�j}=/�Ut�&%��g�]�׺������]�В��?q�s1�@p8����jHDT����m�3��O���7U���N�g����6���[)��v�����>�VR�i����D���7��u1�m�M�:e�(	��b��i�>��${�8��Z&%��U��3)�4bW���9���X�jW���.�TW�ԙ!�pv
�xo��X{���m:�&��{�Eܹ�D����|^k��զX�i+�~�LEfװ�N�OV�z�?�v��;�Gz K���:��^���A�4\'��
s��Z�L�k���wb�$>	3��Z�]���,*��^��&��<u�B��l>� �Lr3��˶���]MT�$B�+�2"�� 2�9ƛz�	~jH,fZv����AK��!��)��ǥ��`������ک0h\�R���
������椝�1G_�p���Ƌc3Mh�� O; F墱����%���Ω�B�S�V�ajwnwl�lk����#�F焿��|�]�����9� 3�Gn�_���Ʉ����r��-7l�*��ڋU� ��[Ț�m8����56���!�LT�(�1ӫ{<C���� y����W>	������
ʛ�38吧(~P�7z"�����iI��������ƚe
çB<J�!
p�Jf� p��3�`K{z�)HaE{�2��y僢~$�4�ͅ[U��`�g�Ӹ���s�*yn�ᴜ�6�kj`6�WBg������^&R,��.��6^ ȱ_T
��	��~i;]\p�XlxVHYEB    fa00     f50��s�
�,�)��צ<�M��!�A��%̏���ɮ�7�Y&2�R
V�R�q����7&����~�E�؁E���\���6,�ٚrw�g(��FyB����k�ʥA''��7�~}��d��'�N}�s4�lˆr��	%���RQHT���I�7د*sp��w�ҽb=<�
��>���I͟٪�.��J��e���Ʉܼ��1��}O��ά�u$l�4!,T��;&cW'	��9[e�+E�dA�T'n�$�߸#޸�2P5�8^�w/��T�ߴ�1�X��c
%@��+ }q��&�K�R ��o6��eI@�_�#�'4=� kZ�b�I��܅�ُ�9TR�:+6M���+��5n��є�iB��� �T_E����F:o�ރ�vu��0�A�:N�@Z�j8̰�����'(E��j�6�t���m_��@ᄺ���H�����4Q�*���2׏b���2mt���g�S�Q�y�Ҹ����;�vb��?���nT�\�w�ż*҆��٪���f >PV{n�W����  ������� lh����h�Z�B�����j�A}k�*�n:r��� U�v���{��CY}U�A�󦣲=Ѕ|�2��x� 8�"�;а�ΗbՃ`�N|M:�D��!gˑ�6�B�]��{�u�m6����o:sR��|�*��\�A�@�2��(WO�%iC�vR]���+pe(�2�/J#��~���śUMNO��K�M3�ב5�۲�x�*)WT8P/�d���]4Vv+��\�Ԁ��{��g]J�R��:�n�1�f*�}��2/�-I��A4� �3���r�����k`n�(��~��)�f+{���B�@������J��-�<���"i0��Q�8[�7͕;Ż#�ţ�LӺ� Df�Q�2]�q�̃Y�\�h)��P������`���S�Jd웞Ϋ�&n�!���W��x5ͣ��C�����mLו�3#֍u���n���ah�(�ȉG�}�����#L~�rm��a�Ž�<05w���5?��<j���H�4˚x�樒~���M����%A�#vǡ��TQ����;&S�o�<��0<P"�\�ו�FB�j�	�"W[\�n9 �U��˾!�1�8/z� �g�^$7���&����bü�G �1�t���/��bl	-Ζ�c��w�&R�v�V��CUU[FCDZ�Rt�g�:�́��K�{Q�	;�@m���N�$��Go?Nٴ�X��������2��]I�������.�$p�����:*�T�T=���Q,�٠�p��0���o�1�IM
9'x3FC:z�n��ܓ�Oq�B'H;E�	�Q xGb���Ukq�йa��?��׉�\.�/ �U}%kc�kJw|KC;<��V��br�5��q�W.+�*����D7?�gHӔ��/�x���.��gv���X:���������%�7��T � ^�_���R�)�% #6��/��	(A�ݞCC�TcR/�d�?���MC'���*M�\f$�>P��I��u�z�Y
��'Ӕ2�x����֝.����8�'���B�*EE@�,���)�㙠���d�U�!��Q�����͢�e :��h$����n/q�mLӐ�]��kj���｜�9?�)�,)�Ŏ�*K��=�zK���P����^����R�%�%�6?P�� #e�~j4�I�3*]�Q�s�.�������:96e��3恅!ְɱ₀y�qw���k���M�����H���X�����/�4}�~����9Pw�F�P�=�[mF7pt� �����$VA'�"��7�?2�o����
7Ն ��=1Q���|ҧ��K��5/�uysJ�._η��]�i�s�b�J^r1�p�������þ��"C��t/�讃���qx�hTr������l]ՄOeb�i2fv��Ȕ9f� ������4V���R�1�0�������eG�d�)H0���X7 ��<�1T󣹝�	�=
��fߐ���_��Qձ2���"{����l�?�eR^0�iBzE��߅�Ǘ�3J���,�HY�5�5����?�`�aa��}ͻ_�����s�T��6YOE�����B�%��)�ظR=��Aаx���HA%!���t#����<�H�^;b! p�R���s�(1�1��e <Uօ�4|O����O4�
P�����vR�)��0$�.O���g^����+�h`�e����h�������a�v�#�kW��y���c�fO�?�sLw�%/�-J��NO)�c�Y�"
{qx��������<��M�?�`�gb���ԓ�.��}�l�0--�l{�Qж��7@^u	����̏��ƌ�bݚ���=�x׍S�-r�b�T�30|�A}95h��&go`)�aǼjL�Ġ}�`��W�K���+�?�io�P��n��S7�vR���@�����g�d�������Q�15G�A\Ϛ�k��R�8����0������_��Ϻ+��s(��-�A(D�a9��Q���u���@�?er�GXFN0��L,�n�ln��l"XF���\��L�mrUV��mN��B�V�������O���ݳ��dX�:��O��uy�Ғ���8`2��6�,?�ނ�i�6�Lpj(i���Lu�p�GU�ɍ�\�ʖ��?�WÁ��Z��#>���]��t��^#��W�)�d�kp�QJ�H_�{�t-A���C���Aq�GK���U"�w�q�+ӑ>�&��2!����2� �'|O�	/�r1��*!d���e��3h'ԑ�� �^���K&�6F��U����4�֕�{��M*�4��:csFm��6���������4XԒ�!��z �wQP��;M���v=��I�zz�]��ڏ��1����D̀'"]��NQ�{��d�\��|�n@p��3O�R"��u�@��%"w��L�r����t�xͻ�Z����`䴝��O�9X4l�!�����룶�E�6���z���,o�-{[ٔ�� 䤇��O�n4��H����4��?�X\sG��Cܺ�s�SM��OF;��hSzOF���ǵ�DP[g�T �y�$�������m��[�t@���q����8J30���j�##�W�m�мr�
%=U� ��̋z�63�]�fqH \I�\�lq\�Ʌ'������y�/)�#�K"/���ܿ��h�R8e��R̰�X���
7��q�tm��g�)��O����6k��0�j#��]������5N��!���t�fn��~�vխ8�OT*)C`^u"���;�b&*���;�LS���_L�y��Jz��e��R�B���K Ș�F+��$�B����)��Z~�6u�W��g(
��@���r�N��8�K�u|�����ܰ�سѬ�ы�VF������O���[1D����
�D|$�z�"������m���t�ҩH��B�T�s�N��[c�c�.� +@�����Ft7���H��@-$���E�� �i���Wr̯��Ive/+
����N�ibt���a��C)�Q��szU��;��6��)x0z�����?~�Q�\���Sw#-�֒��i�  ��H
,�!Eg����K�a`T�z��Ff����|�����.5�-���z%��_� ����гJ;#J@@j9JC�Aas �e�w�j�l����i�}/nC��^��t�l�ch�u�|w�����9��{�e�1D�u�Ŏ�����z�R��!���3I����,�nz0a1����\�;�`A��v���?G/E��?��Uh�+��rv&��F8�j�Ǵ3�3"1���.�XlxVHYEB    7273     560Ww9��f�e�:�\VFI�2O�E�eX,j���s�oc��o�̬��O�C��x��sɖ���b�H�%��ӜA`�#]"W)CmK �S�E����ȋ��iIF�x���ލe��O+� q�#�5>+�9yd��V�G�Y��K-|��YD���g�k~'��|C��w���YLCu�*��kS���![�Q��*����3�_�nOQ��_����-6rq4*����4�I]��{۪��D�s���.mr�ƃ^]S8AFy���&��8���nX��F7/j�����Θx5� =O��8lr��3�/��T�/ ���P�C<������ٛ��9�/>�"YT�=�H�V�� ��}U ^�߰�g 7.�D��3Q�~��;xJڌ��}+rqn���� �m(r廀δ�ڬ��8�Ԝ	��9�f�-��SMV!����hφ�؁h�+FHU��B�/֩�9�Yvw��u,r��7�>jU���k��c45�!���$+0��8��夤?��L/��a�Q��|`˴e�F��Fd�3���4]%
��Xi����A�#�/�9��E��ʖ��D>��6�hX����W�A3�fKti��*���u�s{Q�i�!F��jȁ�33��7�ٸ�����N$�X�9.��d]��z�����Q��J�^��J���a���ۀ*�L�G�+V�0m�X����^��	�{�z���?��%�h�KDH\���p�C#	t�?��� i���0C-�s�R��wʹ��4v>c��Y�� �}|�m��t��mJߋ��y�T�L��q�n}�Ӯ�C�,Wr�`��W�E?���s��T�X��N���k%�q/2� ��C3\p[w��5f��X��S��6��˩Ɨ�Ew��[�%v���&�j��F����4,Yp�AW^��@Z��JP��P[�@d����=����ᛰ�OJd�ꕘp��@BtD�j�IԦ1��B{�:p"��P�`Eb��,��b�=�8$K/�Kc��:�J��{��E�Ŭ��>ɕ���.��NT����v�XʖV�¨�Ӝ�8MՕ����s�L�h��x�v�"�:�����l�Bd�:T9H�x��ʺU�H�t��N�ߺ����6��(n��m�3������ail�dD�F�!�gd'6�\��Gmkm��:뽞�/<3��T.�>��9��?�9��� ����Q�G�P��܀}��� (D�m'�1�ҌS�<�B���	��2�)���`�_�2Sl����g�9��7�D���(��3�T��zR"��k���c�,qɨ�Q�=�Ud۟������n��o�Y�����G1&�ѕM�R