XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^����3p��� B�$r�M��S@T<g�!��c�.ӕ+h�I%Y?��A�9���w�Mu���5�66�L�mN� �h_L�d�HӾ����1	1<3_��:
N��{���f6�U��� ���6�k�g�5��W|�I�׸�R�
����?|��\o6��bj!�'g��ɋ�b}��ɔ���2p�g!o�!=��;�>�.�b*O�:�����ooX|AX,�W�$��*����϶�6V����E1�}1zrY��ɐ��?L�䭼X�Fj�Cʦ�t���0����UWP^3�^_��?�;��ۅ����!����g�[
�Փ|ɲ�|Jӥצ���0	L�/?i�S�Dr�,o.'x��='�e�<-��z�:� �ޖ��� ���oh������F��2ۂ�$�;�{�|�˄�~�+}�hc��f�����#3�t��s_L�)�ƹ��e�Z��%06[�%�bC�5�?���	�U��Y!���)f�i9��G��,�[���xn�)D5�7�M]o�R�n�Y_��?��(8=����3s�|�@c�k��²�*�{�}#N����
FD���F\�#���9Rc#旗W�$Y���$�����,[���d��ыMe� ��Å"�RX9����;G�vk���f,�Q�5¦��9�i�L��<�����#�R&�po����jO%ۼ��¤{E6�xo�� �"�*տ��ڱ��9���U)CςO]r��IiS�Д��,��5ږ��#R��ƒ�ZXlxVHYEB    fa00    1ca0ݐ��$��ߺ9�aIOǹ��y��/_G/�M"�q�_u� ,��Pg�
E[�<�ՙ��@57v� oy	��
�F��S|ݿ��a�����>��k��/�ɧ%�3R�=��ͧUζ�jB�Nj��BG��G���V]�˭DL��-6��,nM"���վ�s��'4b�-�hG� ��{���$����l:3�huA��q�[��n1���.;�D����[���!5/���{�t����������6"��ض�c�#��fE3��ĽR��O |���EX������ȁ�ő�����Z�s�"o�[�W<��������џ�����:�H���҈�V �P��)��9{��wN�b&t�l�I�wԂ(o��@��dU:����h���������RENk�,�*���ȏ��Z�?F�=Q?��6=-���(Ż���T�#h.r���>�G��$��.w�GT}��@B2��o5���j=Wl���.ee�Ќ�8��:�䤯���4^����x�̩̀W{���bUPD���"d8\M6|��������K�,��-���i>$5#�}�����L���g�yO0����4�ݑ��
a��ZL��Jv�
�Q�w�d�ԭ��K����B�������������{�?���%ٚ�m)O<��R_�ߣ���C�3Em��N^V��7^�
�����0���`�u)���
9�����Z&�G��Hꂳ�Xض²{=��� �A�����s
��tF��'���J�[������Q�Ȱy{���$��]��G���u.'>~����Qt����`,0𢆊�i�1�8E&C�h���)�L��4��24��ğ�׸���6p` �_w*	���4�XnVl��<W��A�<�m�7��kj��	y�hyΥ�K���\���O��n��%�^k'��tG�[�~jN�b�
��v���?��McXa�9)R��_���:9�1�/�7��P��o�<���H�z�wN]3 ?oq�7��&Z��U�z���1)+i"$y�e�'��K�E��K��+�4���B�Ċ^l�M�Ò��,���L����V��:�B���+�@D7��W��iH��7�d2�Ae�vZ�~)�@+�Z$�`��ڭ�RѴ� M&� �4�j�澇�~ήF����b�����O��^�
�o��-��2��Y�"W�(�(�=��KJ�\;L� 8x�%������Uj\�w}??$r���d�#�_�Q4�ot;��}�L@�9y�<�n���!]�$/�I�r��7F˳���)�h0��:z�.�bؘ(�7M$�w���{|
}o=��ʁ�ɽ�y�e�d>H��㑗"6�&u
����ڠ��g0{k��p1�p��T���	M�?MY�T��{����?�d'\���﷽������O�&jR3���>�D3��3r����O㒇`>��{��Vr/׉�8	�,èj&5t�dΚ�_ĕvbvbm h�����s��SF��
�2�<0.@}�-�	�}�yp��/�F���P%� ���"�6��n��\g*8�!G�G�@�i����Ͻ�I�ӆ{�L�+W00�SX���N^���K�y��s���q����^��^��`d4$P��.<Y�mxҖ�o���gI�X?DJ��i��4���)U�U��w�1�mq�iJ���ܕ�{�Ȫٳ�1�����>Ў�Cd�iL�z���^�`���	;5v�������aݺ�ս��C�P� _��%��!��ki(�_%�˔�>�)�l
E�-���(B����s �_>�xcW�,�-zM���b�n�U��h�l;~g�0F���E���ь��f��9�����.�B�/�+� ���~�Ë��7пq	�v�����^����Zb�]-�J��Y
M�0�t���5I�)ĬD,�)�ga�� ��u����x���r��W�`H���eUa�=9�e�F)|�v����U��}�-h�\y-7l���2�ђ���)��G�Xv���� ̷�a6�i�ۤ1KF9Y���p�N�'�l���rJ���}?�E0��[�x�9v��߬w7�OZB�'��MG���_��o�t�K���_,���Mt1�`��H��f��_6?��������$|����)�|8�7�CS.Ho��΋�ts,����?�	���K��pD�ʋ�|x����f�pה��1�1o�A�TB�P/I��D�Q1�m[0�������8j�����Gv�@[�X��~q���9�w��t��؁Kwע�̏��
�P-;��IV�/����N3���e΋zK��MJah�ۊ��TB����~�b�?O����S�����P��M��؀�
L��'�r��޶6m'�e��<
5��
 �gd\'�,��/�3ټ�ŞC�mP�4�8ږ��'O�{�9CƍA���ŮG
���Xu1J�Z�2�k$aC�s3���8�r��v�������f�d�g&���9�'`�|���|�f��A\��6*������Y_����3�[�xa�yaֆ�)�n��J����<����/����e(et�N�ȘNRk՟�~�՚[T&�]�BNz!Q�!Lk�]���9[�e�3pA�0<�駑O.n�|�R�UG.H\���ioe�h�eH�m�zF���E���~z\�o����6(�V�&����e �i!�K�H����<� �+V�̹��cK��6E)�=���QkBF�p���H��b}��^}����K8���c�t������1��{�4�|M\g,������˺��G:H��~v���2r�jd��9�?Ly�TJH� �<8���}��O3��Uݲ���"(�S�5�ՌخN��7���G�l��x��۩���,�	���B)In�u����a\2k&�_�o8M�����ng
��&��*�I�a	��G����g�� �xX#��r�[x���u�zǭ�8�������0|^T��� #�0��>"�Dy�i"L�=������4�����oy���N2m���'n�#��u�>>�o2P&��Ǹ�q��'�6�K�ǅ��R�����������:y&�ѻ+3���HTtg�[�IIA������Q�����i�������u�+�c������-A�JRz�w� c���E��Z���r��k.��A��me�4�˗��=MW��dt���{`�7A�gr���y#eCA��VF�A���A�s�^]V�m<<�زL�<������c۴���Y�ۨ.�;�'�>&o4�G�#FCv�9�����"���@�\��Gq�c���)�!�[%�{����d��\�Ϡ��B�QOM�3�;?���E�G�1�|=fD�	֐���d��V�����)0M2��{5N�j��\>�c�N,X�l�zX��ɨh��~�O���>���dnng���rdh�+��T/�eS硅�Aj���LL����XO��Kف�\�'�ǘ&��/��p��ָu@�	�9&�Ѐ��a���6���?&>H�nI��G�` ��+���ު
����O�b�H]�\,_��oXl���� F���#��F��_jW��l���xVD���g�b���Q�I����bk�j�L�h*i�[�X�Ȱ܈VƧp'�!x�h'�&�e��g�j��On
��g�~�%�/�x3�ݴMoT�B��0��.�ɟTt��t"��L�/t�"F�������hBV1��b��E�T��5{a��mJ����,ԡE�,L����^)�����˯D��`�i]/�2߻��ΐ�dsѱ��'�-�����<��C���Y��<7�t�8F���/��Z��w��W�\?I��<�-�+ �k�?0�2�@�)P<J�W�M$�՞,����i7�`L��֊e"0X��^릑��� K�1D�B_�3�v��(�~��nv&<#_CBŒ*��8�3naR�6�5a ��"�d;�|� ��~gx���ZdaQ�thj�ZX��e�T�Ү�ؼ�9��b�[W�G���)��Z��E�Η�q�U��)W��i�E�֤c�k�A�|�8L��&����[R={<\��rW�a�RN  �%c��)�W�M>��]��F�/�6�U��ڛ+/^ð���r�|Л�+۔�
�廼��\)�iF�ZW�;�>�|��LDr���ҁ�ޢ8{He@$W6"`�x����`����#)3�R���m��Sx��q(ֈ@c�����]�NM�A�����Pk�~�$���0��l�Yb��C�3ޮ�� P��)(�s��+���G������&m��T�M��|S��姝�3�W� f�Ƌ�*}\N�,pu*��}|/qٿ���Y������A�4���\�B�'w��n�=i;�rQ45�+�S����3��2�2�6r�kWT�Pk��G<e��`�����Ӊ�l�%TEZ$5�&K�[�P�Qa����Ƀ���� ,��$����b�?�<��8<5�t"���!�À��#�J��Z�\[��::��j��fX����=�t��ؘ�������؇�i���UW�����s���;�i��仺W4�_҉��}��;'�a�#M؊�*<A��:�|����(=��ˌj��	P��/S�S�@����P<R�K�锭?�5��ay���%����#wk}]�n@�=!2X�қ�[0�{*	��)���F�@�)�E�S�m�7� f6�+]IbD�=�q}��9A�=tW��T��^S[�zͅFbܺ�)���GWCq�Q�VAҝ�r��Zo�@���u`zWᨚ~;�����O ��z�m��W��KXo)��r�quJ���\Z�Q��m_D��M���J�^s�g���	������T�+W��jV
9|b��Wh巯���C�x��9`����Bj+����?t��W�%���4�i���hH�����\�]�0��w��"޽�]gOj��[=
�:�J\�ҟ����@mHst)��4#�ӖKP$�@�r�ֿ?@d1���Ie�.����1�Z������Z�xs#�A[ZT��L���X?ذ�헤� 8,�ߡ{E�L]�C�~�Ad�����lVL�,���f\�=�,��/Nʿ;ojT�rx����S�,�ev��}or��5������&'�.v{�X�l�Sz�Bֽ�Z��u+�p�\\a[���rȇ���2��Dߒb?&b`������D�p�6���P9٘�,��S)
�4F� &�b���� �٠�`ъ(��"X��;0N�ޚ�����t�żӳj�|�˳YSXVa�ϸm=�?_h"*|�⺏v���g��R��w��jm��@�PM���pKmg��d�l���ut]�<�0�|���&G4���5��cTL�z�m߃�D�@P_\���i�.�1��2u�P֏��˰y&�b���֮��s�M��Smq��`���"�Z��!�%R�	�:�>ꢛ�����FIC-yh��
RE;�Rw��y��?J�M�4��a���YL5���d(yg�(ƉN��߶��F�Gl&��]�����6S�-ϗ�<��7H	�S���)�GT6��9��O��]���׌����wz?�x����]���Xa�Xlkh�:��-`���X�JJ����Z�����Wf��VWH�������v�H�}H
%��:t��vɥß�C�A��y�D�۠�	��x|��/�'<�ZM�ۀ�ۙȿWI�N۰����Z�X��G����8ir�{�P�oB�r����W�p{x����,`$��N��
�,j�bGLy������tAb�k���Zb��z��U���c���B^�g�q��w1��!����[嬫��N)
t >C�� fM�)� '`�-JI����W=qI����m�~\nz�FHj�mp�{!:���(��oLr:_&�5C���Y/ussc�%Ro����,+Z������5��~\԰{�h|1����Rr��8V�)@"z���<S�؊�F��Z�������CZF]��{��j"�g�����?��<};js�B ��js]Z[O�1���ucE�X���1��g�4�3dh�Z.�����C�E�#�J %�D�1�,m�VnàZ�4��5��0:Al^C	*v��u�������Q��&�7\]�H�R����ʩ[Y��l�ס�%�� Df�2�k�@{y��M�Qz���!�;Q�
uRc��S�a;l�)���3�]:�gGC��4��(?W�1֬ꘘ��P��Df!�jX�bj�&�����z�'�o]U�RQ!��rl�K�i�/����tqRW��I����Yno��8⹔9�aJ
�&�As�6�Ч\9� v�u�?�_Mg|��Ez���^�|XiUl@� eS�nw]w2����n�v��{߰���~����x�Ϻ����bj=hc��H��z����SʘX�$&]� ʺ�	'V�Ol$�QF@9��4�B�J5rL�R��Y����8lh�>�P��D������#���\p#�ǥ8\v-��ca�I#�?���[ K�B		��B���T��ŉ�) [�>����H���DA�\j!c'rmY��N &'U�'Q�p�^���1-~���9$i���PR�t����K���OՅnHѸ7��2��6�-g%�y��IM���M�¦1l�'���x�����Kc�֐J�"e� ���N>�۞�c�l���u���c^&�������u�nF��kH��`ažK/���en�T<�A�d,k46��#N`�$�$�R(�l)�j�r��{XɆ�x!B�5�`�[����z|�P ���4�*g��ር0ԾZEfH8�bm�~��Ow-�)�|{J�ܺ�,�l�]�SM��!� ��k�4����|���nч�S�?�Yp�����Q��V����.Ɠ��e�_Rꔠ��;+�@��,�!{]��Eyo����� ���l%���J�Q��I�]�C���"K��н�h�/���uD"�Sp+�nd0
d�o��D��:t!�\c�{��=�-��Ѥ��(�Ie�V8����g#U&SP{#*'�k)�<�ш&(+m猋fEw�@��=�6l_��}��&��Kƒv�쒔����U0فľQ�F�"T�=������W8)�.�K��88�)p$�>���<>�;����j�z}Om�Wd�����|{ap��)���D{�P��MC��XlxVHYEB    fa00     cf0'4Oy�F�
��U��^�\�H�ؗo{��>� )������au��k�?���2ȇ�jU�
m|��Ƀ�(����Ӭ�;��{�
`���e߬HT=�:��`jx�w������� ��0�O��3�ƞfU����V�hB�G�r���E��d�A���S��m3�@x�#�}��<�vd��1'8=�"�`%am��1SRm[<�pЀa���h����1U��P^��K����~��b�oW�	6e��K*\P/���t'o��R���J�ì���`9����&b����x���M�6��F�@^�@����wآ��D�=�ҭ��g�c
� �J(����$�V!~��ƣ�3p��.<Y����5O��4���M�/�3am=�	.w�֍D�I,���#��݌Ѓr:�t�.��D*�ϓ�K I��/��l���%0?>sf�)�b۝��BY�c�"������K����߼�z��8�T%\o���-��Ǧ=�K!�����J��`�ش#��y�!c ��GH#T��i�թ�K�١�*��H�{Kw��u*�I�a�~4�Y�׭)y��<V��V�I���[X=N�-X����4XN"N�鮹��B��׏��=ڑ��C;��>�jI���n\���y���5if2�%�M����uX%���~�LpٽE�B��Z�S��:��Ӌ�ELV'L���2c�|-��P�}�[�D'��mx�fl��D�ޤW��1��k_"�>Z6j_����n,U[��g(R��(°� �����uu�'�P"��۫^'S��LG�3�SR�!X�C�)�D���� ���su�m@:	�>��|��3,���4���W[�9삊k�?a>[�4�H�.wr�^E��X6g�÷?�&�^_T�Τ���b��̥@|�׷����?5��7��R�b������0e�A���bS"M%@9ӟ�uC�}��W?!�}*�%��%9�)3�����%U���vD�&����#�'`F>YP�rQz��Y�6,�`��S�x}�3��+,�uM���/��O��}���y����6j�W���<���s�O#guNL�Ɣu�;=
�A8gL7Ĭ[̃�H�Fʪ����C;G�zӌ���F}�z��ü���&��Ca�"��F;��>_�=��",��F�y_���Opm�P2h���O�Fg����
���73��t��	|>�p�.��H1+�����M���p�t�d�<ܲ��S��J���d�eח�����n&��D�{���qP܁q1����p��A#-Ce��@e[qͪ�K�O�&*�h!��"tb����`�Yʧ��<�N�9
ϯ�OХ&���o�TF���u�A��@�of�!_���Ԁ�j`igK�`O/4g�^�@E�0��QP�:�m���]1)�{|rc�D�Y��'�
�/̱{\d��N�.�`}p�p#7}�(V�'�o5v�J_��hLbk�8�e՗L;&%}V����v=���1����t�{�jf�}���E≏L�I)(�>�e�+�C�]�R�f�1f����b��c�LVMA�1o�8��P"�8O���~�_�[Β��G����lVS��f?r�k�e�Nzʹ��p�O����D�-}���,ػ�v$�]h�	L k�S���}Q/j�m���7_|iā�u���R^l�/��h��ß�k�@���.n�����~L-]gЇ��g��=����ZX?��Pj�.�6�C ��M������$���x(���5����������_�5�=�۵�������$�A<�����uY3k*�iK�O�����$0���x��^P���Aw�{��s�L�����UL�٥<���"0��ҭ�$���3��4����Yy��W�����\'|���6�,�2b��k.�O2�VP����4����[��њ�'A�P0�ʮ�s~vx{_>�E��S	���k/p��q;M.�8��Ja<�������_�O�nƿ��:��y���zu*k�[�<Zu/�U�Z��L�G}��vƃl��xh�N��+a�<���jaKE�>�>]=�{rOqs\�Se+����V��G�~�[RG*X���I����0AHxT9�(�a���%�N�����vNYO-C?b}���7�c�y޹J���Z��$"�!U�F"lM��@O���" �Bg"������
a��#�T�L]����*7�.��d|@m��֑�յ�K�N���57q9b�I����k��t� ����rf�onW�~�Z%]�Mm�朗Ҳ��-�A���(?�%�R�����;��'��R�z�˻m	�ץ޿:6�����wQ����.!73�p��Y-0���/�|TRO�>�GO�X���E����e�UM��>lS\�1�6��J�O�W�U�PT���^N�?Q]��f	3C3�Ve�>ҼW�}l/R����ylQ�zrA~3�����,�n�n�t~��+�k��4��\k��O��vI.}na��d��1���䳐o{���Rh�bZ�S2�s���-P.���0����g�1�2Һk�ɡ�,ή�/f;s�
��V��	5�^v�e����$�������'�H��3"�A�w�`�w0��_�$*�G��"m��a^dѯ��lDd����v&z�6�j�@ O��l���;b`�$9
��n�x��"���OF�!I�<����<�SӘ�W$M	��8>�s��D�;*{��aG|��CU� bd�������ՉfL��UM���09X�W=�[�:��:&��S����-	G���oN�my��`ϏEL���g߳���K��>]�a��t��x{�cOſ�]��j7�2S���=�K�/}�&2�=��"(�b[`���\Q	ޜ�ո�H��I'��Ĕ2�9	@�S3�~�T0q�N��
��m7����<>����V���o�L��Q��3:�i�#��B���2����T��
��kT,$�wz��[�983����$+T�_tD��P�ػ/��&ЗM7�Mt���
�����pk+�'��\ؒ�j�߳�!qf���Ɛ&K�g�}d�I�d�s�G����B�6�w(���HWC���Ho�-3�U�w��xa�.�CJ�����bض�d�xf�"�Iiy�؊� �Ph@�h�����%7//����r���XY3	�wF��f���r��
|4�QM!��P�8:��S;��ܓ��@�*�"/����G�ƫz�&IC )1�2ͺ���W��TJ@L��T�XlxVHYEB    3981     4d0���Rr@�-�P�C�|}p�~��\���g?��BV�x�Y*x��36�QA�v�9���ĥ?�������&4��[V�Z��L<W�����������e+iƖ��C�h��wu������)xI��ซ76�Ӕ����(�����Nr��x��^7/jWP����T��T����86�ͯ�P���{L-��ȷ)#A�Ѓ?�y���
��?h/���y��ò7���h�!.�ru�����L,3??�4^��a6�}�P����7��b�G{£s��m��z � %^?�!4�N��>�+�(�Jǒ�O�
C��j���
�c�+��ބ7׹���.�����v�kj�nhӠ�g��������Ex=?mۅ&�Y!��r�)l�6��`�u>(�y�z���i���R���aPn����nP��7W�����n��d���E��"(���w�oc	��(3��:��g�8ۇ^)�߭����a]�X�
�Y�B��h�jËg��Y�W ��9}�� �9V�C_4��>ݬ���l��H|�EO~nC�ǭ�!(��f���1!�b����8��/�_)]o�?
ԣ�����(�+���1��mۗ��@��j)L/]!uXg�=	�Gھ͚�k�n�7��t�Z[,�$U�_}֋�F��6G���7�ò���r=���(���9j���b���: ��dfRi�A��Cժm��:��gz5+JKdB�w��j<9�h�σ����9AYgXTH�h�mD���z�0��M@a���x�s�1�K&(�za����G�q`�^�a�����u����z�M�'�� ��r���2z�7�ŨA�fĄ�<� �,���&����Ƭ�{8gp�.�L�I�S2E@e)P�}[����p������z���84d��eub��/�%m��	٣��w�]���Ƥv��
o�!���9{�I��M�I�2��+�̰i��<��H�|�
���t�}�H�|5�{y7�Zs����\�����d"7�P8)U�g+����V�g��5��3J�A��S�Ai0�y�c��Qu��*) ����oaz�������1��U2���3�ȹ�X��)o1蹣�ý�����96z���=�ٍ�W2�5i�����B��D���9 sd�|BmFٜ_���U-kz���s��!//�<�X�J��/,ZX�_yQ�M