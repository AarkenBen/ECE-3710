XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3e�GG�͵��y9�E�G�(�t34|��E����]t9@��K�2�+���g{Ci��Ҋ~XL+��R����>ti���`��l1��k�@-Ry��9��gb*;�v/Mo�+�`0�� ����TC4$�9��0��H��+h'����
���}�� �}���|Ӊ�U��:Z� BT�oHF��(ܐKi�2]�+�q�s{��3D{Ư�*�3�! �;��ރ�6����8$�	9*�PE�e�ihr䄟�4���ΜnG�����b���c��P���e�L�)&).A%�}yә�Y}���c��w_:��6d:=j ��u��JZy�f��է��j+-AY/u���iۧ]�0����I�^�աO���&�r��������z��~���D�F吪��-s�����>��f㛔��K�4\~	I�a�
c�3�哀�	F��7dyRɊ�µ�G?H�j��)_�����M��R��w�q���H��0���q��*���n����%@���׾I���m��l5[���vi�w �|�~���z=��Q���	����Z���g�i&��<̽� kU�<�N����ƚ���HW+
�R���E�<�ђ��0��|���h��L��S�"G*QT�n�*�ON(4
��3�gہ�����N�- �z�\0^�u��ڌ��'��G����ˌa�Ý~2�qֻ�Q<z�)��FL�{�C��j!��wΊ��M1f��e1�&e�-�]Ï������l_XlxVHYEB    fa00    2470	��|"݇�Q�ѕ_��3��5?�g3=�w���Z �ˢ*X��b��kl�=��7C;�I}�]r`����2 ����B��}�+�Q�c��`�q����?�0���!���u�ǰA+��l���(��P�4� ���C�@ ��B�>��j���CLqع"'C����*��ǴkiA�hd���"��;hc��s�Cm=)Z�g�q˗d����9ɤ����tqFcQ��GD�qR��s�Q����È�#e���3�.��vY���_���#ׁ��{�uoK�2��Soώ=��B5�t�������� ��\��m�A_0���s��4���� �ÔYH� c�}�;D&��͘6�N�K4YzNFm*�k��Xgm{�:6&���j�i^��"������ύ�}⵪J"���/�\fx���"ב�b�D^��|+���d7g�Պ�߳�gC:Kx������x�;�=�"K��ߋ��7�\�ɦ^�����J�.Ѩ.cA�<e+1С��0���sEK�;3� ��k+~�Ӕ8k��r0�6u��L���Z��Gc�,ϡר��,�*�#�'~��1�X U����nLa�g���
�|�l��;y.�]v8��jl�|����/�Ո���;����A8�L~��x�n>ϊ�(�z:�;!�Tfh����:��pڏ��v�@�:����;}�=���կGƥ��a.N1Д�(�!�nFؿ�;�}�;ͩ�5���8�par'[��P����Bp���G��u �--�:S���nԪ��sY�ќ��/���T c�#��[!����I�����Df�Rb5�M&��@���	:i�m�kE�)������L��`Y��k6Zڲ�\�
'2&Ա�ӯ7�ڤܰ�g�WT��ka%�?h���m�>�[���s�K<�2O�E�h���}=��"g�?����]eǐ{��u�i>H8��P���A� �c�Y
��*������_��6�Ŗ[���j���V�2?��2�F����y�pѨ5���|��.�ؔ�ԷG?Y󸾱��M����;�ďQ8�Ǒ���ogdj4��E\�-rͲ`P2����ږɶ����TaKď����7 FG3����O��d$>�Ӈ������=����g#�U·�ָ���PU�R��ۦM��F����]n]8F	�P�C	ޅ4�QK�s�sO��i�1z��ibL�CM�F-� l"���g���I�0l%��o��b�'�#i	)�9�E�T����f�B���Վ���M�/O�~�A�&��~y(ٖ��L55�M�Y��$�aY�f8t��0�!/h��^e �n�vL,P��^a��a��W��ĉQ�����%�P��$��zd㵶V!J �gbK*8__��;:pw�� �V[�<ӟ|P~�!	G5QJ�.%k�&�j��W�Z_�AE0�ޥs~���N�[�UU� ѽ!�-�@��b��L��m������3D���i�n��l��"���ھ��Y��N�d�x�z'�U���B6Gw[9ezvZ��qJg]@N^O�c��X��U�;Ɋ¹HZ?jTík	1��&%U�������Q�溱w;"G�l��6�I�k�4��̴�K��l�0��U���Z�mǓ,���d�1�]�}Ư|��'�ֹ�D����y M圍�Ԙ��x��E���)�u�zw� H��������BV�J�����6�g���2$��ՄM]��Ԅ �Ҕh��F�Q����GH��bsiz�R�#S:����[�.kd��Tx�l��j��U`s	���~�؁���t���=g/N��\�(��A�m�r�S`�3d�s���uk���vχ ���FD���Y��B�K������e�c���ԘS���\����E��J�.TtIP3bfD1+hn�	_��U�^�-�t|u^�9�<)x�6�A�1�����d8d������X������.{���AQ�`�U��UEv{1�{���9��f��35Z.ٍ��o-�U��@\b%��4)��� KE!qM�G [�35וK�@s�cs���7,������(��]/�װ~���p�b�^;`�^�O�Ԯ�N���5�<"�{�Y�j\�z�&�l8�똻Y�+�qo\�r&S]<�v�Q�4۶	�6g���&)�˿T��*�� n:<�[?�&ul�� 'ɗiǔ�X�ğ�t ��)"�f��*�����_qoJq��n[��+O6��ؿI,w}��n�i�:aR�}�{�%�d-,D�s�A*����~@�'��_2��� W\Cq��dZ�p�D}TԮd(�� ����t��g�����]�VrQ�=֒��K\F~��k��;`���f������3����I�뢅7#*\g~�H)-CRA���T�g�\�צ�|5�L#�q�����arJy�eJ^V�I����.��z�p��&��-�MVH\^~�"@�Ƥ�X>�p6iŵ?�`�� @�6��?�S�: l��i�ڿu������N�$�_�_2Y�|_Ex�ڃ3���T��%P��qCk"�h+�/�k���i8�F�f���*�D�u!>Į(C�&�e���fhy*
�F��b	LF9��&w�0Z{���_0����pH4O�)�eq{~�=��Yu�6)��J�ƭ Ҳ�V� '�,�����VB��xU�&��jj�A���%�;�����[g�����66�[���@�L�kj��X����qi��,��J9��:�6Q�:,c�S�~�0���_�(�䴭Q�̌JK�(���k��
]��@�6�'�>L���K̆��gXs�Ŝ�uc���|$lAk7�p�B�v�Y��x�~�iߟ�,tB���w��`�I8��0��4��!��g���ѻ+�, hL���ɖ��"w�-����Nd󉍥H^��W�L�Y��� �����c�Y�ζ��8�=4�`DCH�*��8V��m6N¶6PdTt�S +w�|1�W��.'������#N�@g$M���9 �b2���&�0Yg���8!#���A��`H*�BWt������y9��3��[�X��l�B�������w]�I����[�&Ck`�21Arݭ��!/�~��b��C������c��QO�g�����zZY�5)'D�k"|�:��@��{;z_�c�'�i>�Ԉ� ȶ"d�w}>�����F���o&����Ԁ��17��&�u0{U.�9�X�xJAP��ѹ��':9Α��\�V+7���:2�Y�	�
���䣺��	Y�=eVp�Yv�����Þ�ژ�}9*>GDTi�[�i0����{��_��,���9u���UL������=𭁈V�P���H�e1���-HF9� pe���L3";L?�`TF�ξ�|�rO|���Y�{���9�@��D������/�[P1�+��?RU͵����� e�1�W�z��ɑ]�qQ�D�5���'1�93�kک(7�0&�1r�Qo���N�+
8��?�B0�AX��P$%;�fbY�i�Ė�]�K���t/���e8�a��s'���������o�H\R�8��� ��<����`gDp1G@Ĥ����)c�s"n:��M����5�s��'���T<��P��d.7^�,�f2Jq>�g�I��7wT����0S��(��o�,1)e'�����l��i(2��6Wp�ـ�yT��H�ړ4˅���l�TW���|�"x���E�(��Gi�#c�����xAPͤ1|�au-��+l�#J9���C����;,H/k��vu#.���)�s��9��m\>����-t�E&�x�/�'VK��V�����P(d���/�"г�x4�h�b�J1�?zxs{��p(q��ب5f�:H�!���݇ ��ĕ����g[6�3r� ���=W�c��JF��4s'�z�9�x�#�M��'�I�%����8I|����f�Kɀ�DA��1-|U�u7�<i���S�L���M�a�n͐�_X�_��Q� ��h w�y�/Haa]���� &ܦe;������mN����"���Iqg���ˏ�����x7Y��u�a`�O|�!%P����尤����|�Y��}U��5���^D!����T�G�g8*z�U^a���]cf�1#I�Aؕ;��O�PMq@+��:�R���<!�w��\gv��d|�J�S��A�q\���!��Q;��q�O�)��/}��KiF��x���N�Ȩ,�9��!�������R��AD���6m#�6�fl�"6����bYBET`�>3���)\�I�����gp�;�-*.�6��>K~�ՠ�Z���tq���{t� Mw"�X?�����!C�똟����^|-�Zh��x�3��9�԰�-�BN1O,�p�:���C>ʑ�C̅ .���¬F3NP�I-�aB�n��������_�q�⺢��d�ȓM�Jp}�HcqhSH���p �߀���]l�$'��?H����#�F�fH/C}���C���nq<��9V;�Ɂ����y�͹�L�[lޟc�pq���Զ�b�3��h���;�~�}���,�Q�bO�4c�T�|?��;������AcͿk�Rx��V��9�-��ye:��$zIg��r���fRe+�O�c�|`�.�c�sBrhk�~m+TR"��}em�<�$WC�����(a�ԩ��W�ETF�ܜMȑ�%�͸K8U͡oHJ,�>Gk� kc�A�J0nl�>��+�B/�n֯�C��mah�C�9�-�tw߸dE��n+9xc�M��c��r��_u+�6WK�C���C��:%��t	���	׫-�\3�E9��r��4�	"fښ��3X���p�!�M�5y`md��Z���O�-�S�}UG�]&��u�a�^l��o�Ͳqj{N)�-�W76ǂ�T����� ��DO{�Y��*5�:y6W�L�͐�Ł|Ԝy��>��D9����V�� "�#$	�q�Qz�nU��%�g��E��.�VbS�֙�ے�$�<A������P$���&�RY�p�,`c�hB����cO�Ķ�48 rlN�&�����4O�� ���^��e�L��5��������EF$���=�9e4.�
�k�'�=�%��[��qR�Vq�`2yϊL�zg�Wq�?vO>Sa�?�r�9�I�n�rL��p�6�9L�pϡ!�tF1�x�������0���,�ۋQM�n���
�tܶ���hu�ҷ/z������@�p�(��q�(��뺱�	D��	Ik�8||t�^���>CW�S���O���}\wB�L�`�X�&�A���9e�nq���^k�E��H�٭U=���	�֔�lmRĭ�?��z�3ryQH�I��áBW� $�gjR�U���5TC���u���a�B��;C���N8ȏ�	|~۴Ǚ)>Ҹ�AMx�hL���@x1S��׹Ӈ ���3ħ��lrh�����������9��VFՅĒ�}�2�Y�g�-�e��/>���ICU��A�	|fƾX�8$\Xg=A�{�w+�\C�ş�;�F���_W�#���̖�]�QU}�mpO��gX�X����f�dG[��q%��y��e�^)F������V����R�<���y�Z�9��ހL���j�jU� iGA��Ź���M��C�Eԛ�X͡�[���__#��en��h�jg�z�h�a��v�({NJD�������.�ZL�ÐXppZϲ;��q�uj�����7�s9��ೀ�p�aWȧ�@wT�>
Оz��=��S ��.�� E���Z��y�ń������R��:�5������L#bhF�f��CDo�����'_�R�'�; �WqAH��g�t��zF����?0�4��`<�}_;Q2*�\�����|�쩜'N���h�����P�J�Ԍ��Aԑ ���~�TT�Z� ��/$h���X�Z}�������&j��C�V������-
���h�A��/8L�f�޸}�NW�C��S�*Vַ;|؁��
H�N��$��p�#5QEQyʺ?�'Y��IG��|`DjA������: �rHQw��4��J��m����Te��������^<�j\W��'i��i�3;e�!�����/<�˛d뇏HH�u�y�MN���}��5S�ܯ��,�:1���puj��	U@�>�57��  Y��.���\)������$w��������|ݯ�O՘q�aNlf�/��):�M}:��� <RE_s�H��C{�r*)%���ژ��e�ꄖx:�/ƳDk�rEi)rFS>�)+���t���GVZ����,4��?���-�� 2É�)���>є��Iج���J?|�`Tr8�ނ�n�I�=�xÆ�DC Z���z�ƟD6:���-n�C�LN��[ی���­9nqq��;9����yq���b��!����s�����a@�aF/���0a(��2�N~%I�?�N��5\�����d��ҵ6��cW.��,�O�1�(Ya��c��������3��N�vtޘLo5�@)��&gQ( ��߈;:��5���IA�s[���'��ƻ�Oybò��ב�W��<<|�g��q��{]E�ַ �X3J��oޥU�+CN4l#��vO��3%��Ar�ɹ�V�Uw�оp5� G��7uG�c��k��iGe��:xf��@pk�pn4�;�`֖����@�)P���Y�������׋/�;Z֍���	O�7_s�~jA]S�|��~43�a<	���p��;2�b��_vM(<K�.�]3˙��uܥ��^O�@4oq#nb9֧{�a��4� �����K�LaE�[��O&,/p��&м�DV�9�Y��-���&5◐��+���8;�K���=���l֌%��jI�3�^q��{����\�c'��f�UH�覨%l`�\��̡P<#�eDBf?E^ގ ��B��T��.�i��7"�X�R���6�?��ͯ��i�~� 7���ü@k����y�$��V�V.p��nFu�#�u*Z:��i�K2��b�`j�� 7�A�~Y����%5Nbsz��2>d�´�>���p..rXf��F���VUU�WN�|_]1%@�k��B1�$})V�YB@��'��}cC%MNlfŮ�7�G�c�gk�w0~�Ġ|�����SW���Q� �u��$pK'�#G�>����ʶGTV]ӎ���<әDG��ƀ0�?0�|w6� }�����0���Ʀ@�dI��Ԉ,���FU����C\���.I3gxe繸J�׈�PUV��~������)Zl�XP\Ѻ�^'�d�/���A���9���K��8��c�"��Q(<f��EY=��^곸�A�k��R�:���f!��,4Nˀ�Ӑ�����u}����.���RR?��:�
pM2ysƱ��0?e6#¼��_\�<� ��ccTx(�6��e�����B���5�U�g�%Od^�>�$��_+Ω�<�W.�Z3����^�2�"�rܲ��ܗ#�"�|�����hY$����O�� 	�BC>� ��pp�����w�+���Ѵ��Qq���*����S��_��K�����x��p����ݾ�WЛ�VP]i\��*Z�� �#~�����@�ַ�9�9�n<<m��n�a�js�������n=�4mh%��J�5��W�Ŭ[l6�ٺ��w!)�i*���3  �����}lV�_��R=�BJf_#�uȔu�$�d����~:��D����e�6%n�i�����jv��H]H�%�� >v��8+:>�U@�')f/S�T�|z*�ϻ?�5R�3KW��ޭ?X�:U���-�P��O�p>J,g���B%0�u����:��T�����&��]���Y���u82�CB۾��C"�����x�z�%LkD��p����Ru��� 8�Л&~�
�
�L���+Z8}��ڋ9��3�i�m(��]ٕ�A`|��Xs���B���/5NL'�_�o3 |�T�Z��nMc��]��]���֚�f%�n#��%$X��8���|�\X׉W�َM������������!��"���)�e��9�O��f1��kV)�u��D�Λ,A� ��[d���@��	� '5-P���������y�Q�@��-����h�˃����")�}Z:�	�l�j�ᒮ��x�՜���(�������;y�O!�d�Є�
f{�t$q�kr�|�b����Wf�1�lO��M��AD�9��y%��/�����?'�ԉ�h�	�cJ��ow��"�ȳ���z�����O�55J��̯�o3n�Y�>H>�z4�&��e#g�K�1}�_�]<�E��v�)U���x��:OtY�`����ꧦ�~7J'�!G-}��m]vx}`�l;�W�L�v#>Ϯ,��"��Sd�I����N�K3vu���D+���Ċ������;�j��1�BLb�;n4��F��hAs�ک����kA��"o��K�k���ٶ����ł�3>����4�UxN���zM�v��Kw��ʄ��o�7xS ���p~�s5�ز�SUL��d`_-ֲ]g�-��N�����*�A�Zz�4��c��}��XK���H4xj�U�[X7_sf�*����4S��G�rY�]VS|^
�H�+;2���`�K��~߫@B
����-�)��?))�R$P�C�;4�_�dd,^����'��ð,L卋��6~�x�Z��+��a,FLbvRј�1��Z��� �0��I�~d�'{Rm��}2�8�5S,��A������0Oz�^*=����W��!M�d1��f(�{��h%Αs~�LNFp��"AwT9}�e%gM�_s��S|���/�Zj�2���-��-"i,�7.��ϦΘ;�1q�:)���೏/v�D�h�D�d�ؿ-����&OU��ϜϑK�b�3~�L���pS���]DQ��Ҳ�e5�C�Ł�0S΅�:9At��U<P~��H��R	ef{|�IKC7�y$&b��EV�Wp�Q%�٭F�n��	�F
�FS��i��{w"��u<�����,1�߁���Mj����N
A,��SN�#f?�+M�ҺOȋ�9��_Q�9��O�X�Fh|����	V&x�+d�ǋ���gr�X�UGlb+\ɞ��1�1�w!S��Kt�������p��0K����XlxVHYEB    fa00    1b30��d"���L` v�>��/��MB�����ˉ����sZ�"���o�%*e�fi/X�Ye$%�.�&Xm�� c�ԎPQ�<��Ϝ(�ۧ鞈�4����!A�"ʺ��*�sL㰃��N;u��=���I{�B�&D�!_����1w��\��Ȉ�c��S��k6L oᡠ�[�8����i�'�;��Z����� �;/�׼1��G���|b��0���ٱR�~�;4�����301g�b�� #�s ��(̂��~�P�o���L1��W��G���Uܩ\�Yl�)O��-jON���NCp���/���)���};ʅ��.�c�ߗt�	�A���CI��",�s<r!�ͣt.���x��*���Bx-4}=��p�RKd�ʲ� �'7�U1V��}���,�s��7��[�������~��\%3K��;4�!S;yu�U��@K^*Y����%��W�^�̲���WG�#�Lc��>�H�1?�ԉ3;z��p�"��g��n@O���ʡN~!m�<s3����ld��	�ǰ��H�.Bp��'�<�s��g�;�&8Q���y:=���v�Vݛ?����Ѳ^t�����N��߳2��V��:�.u6���xQE�y�kC����E̶���f:��qp��2Q�Nㄒ���}��P�����S]o���Ia٪D��]�^�lB��ܻ:nb̗��|Q��U�B���� ���W�wO���ޝ������J�ب�|	?��ؕ^���^��2z�v`�jZ�]ws'�i�����eˡ�+�y�6���ZG��vg��˼㶥P�%랚�}]��=i�g Qrio��/4,H� �Pʈ�=ܡ��2�p����Bj���<ۃ��#O�<���<��҅�S���ʒa}�P�F�����? d�9�䑟�
�g�}K&�*J0�/�J<�$�g��;U����44Z3���d�˚;�\bkK��AdAr!5��Q��Ɣ	���̯���t�e"w��x.L�	<ڹ�T��R��W�N���X>�Sb4�8��iA�T�6���#�l�|��Ky{�/H�o�1���sP��˷jr̯K�j[�f�������H������;θ_{K�֫�OhaS�'�0γ�|�h����(�+�+VM;Tb&�����Ќ=���$��B��-��ڢ&�Rg���尰�y��lGG_)}(��� -�qò+@�dF���aٛgV]+��?�7��sJ�L)JW�no_�~kd׎�_R�N�I��>\? �
���!�����F��|am�S�J��dRu!�!=1�%{-�tH���ޏ��z�V�O���T�o�m�DfO6�)(�:'��:�BN���?|�]O"�':Hv�f���|�������h	ζ�$_Ѡ�˃�)��\��!Y�e�z�Q[������1��õ���GB��gH�/Je�aH�H�·q�Ƴ�$c7�uʝ��6GO�H�2z�.���-²H���eJ�K�PW�`:m�f�咞�\�4�O��|����y�Ge��uյm4Kc�I��sw�Eb��;��@Sb�Xq��hs��
�F��1B�X��3�Uq't'	�����S�; BOD�FD���DW������tDw�Q���UP��V�����&�هh�J���͛�I-�x_pdU���Ĭj��*y�OբtsB(IH
�p����p3V$c9��}��'x�	(u�T�!����c���|��qw(�S�q��=��Μ�e�WXV��誟9��^ŋ�����ǚ�u�	���$���kt������XAX����T-r�Q�{S�p�No@`.)���.I�>[��oŉ>�E:3<����,g#;ic߀:$7��ܟ��5�j�S����}J�Z��C�я��5l�nٱ�[Ҋ<[��Ց�K���t��
�oɽ����~
d���Spθ�s�$x�=��M���Z���C^�]�h]*Ŕ�ħyD@��v��)���I���u����F��3�|W�ٞ�D�@�=�m����C:9���bo/�&������x
��Av�F�j W[�Ж���fT�qX���-mg�+#����h\�TI�����xM��We{�ȟ>9����* ��<��/�%���w�}y�z2�7�k���gW��q�j#�4��Q\;�b�M�,��C����n?��v��uUL��!?$��'*T�6��c�
Y���o$[b����z���l�������t9�� �ԐJ��'�bi�F��t����Y4ͥ�S��򂌀��]}�����K\2!���8��+�D"�uʺ^��Օ���Y�;i���N�Zn�XM׀N��E݆gR0�������p�iw�����f6�֢/�)�BD"�����cB�����9�.�H"��S,��k3�#J��)���1�D�2~{��uAN������h�<�'�O��42�wBm��<�g�Wd��<x�����DO�5�'��µ��Zr�N�R�sƞ|�gHl"�
I��z��6�1�zM3�e֗�T&��/��>R�6�B��Cg��ӛNh��=��ӛ�`�/�س�~�a:W��Ă��LY�JR<M ,�_Fۍ�� ��jM�U�Ǯ��V'y��j�tM�)<�uA;ܐ���Ե��z[n���`�9�&���.G���u���AM�,|:*�7? Cϱ7_����`V��G��D���B4��t��Z}��H%&�k���+�����Cg���:��\nHa.~�a�����)��*����Q��2��D�&2���<�g�l(5���3�x�xj�v+T��Z>�䔽@��6�p0m(�<���D�/��{<��7��v@̭/��׳�;xg{'�q���E(���U3S�}Ӧ��|�s�W��D�~������+���-Z�����LF��aF&��S���'�,����bCk�ny�kZm���B��J�󃣜ہ<��A68�|�	3˜4��{]=��/��
�Ud���-ޫ�V����oq����b�B��<jc��;T6:P9�K7��z��Ne��(��u6݊���B|��?
��T��C`���,�����N���AEn�E�<��[�K�\A?����U.%�E(&`�gټ�1T��%Ӕu@|H�N8�ޢ�cF]�7Aw��E���g?�9���>��*�.��X��j˦�bW�t@���[x��\�������J��w�`�^3e�#�{�1C8Uz΁��㵋�t�7�ņC	�����-V����`��K,��vx�C�h�܎���7fL�_�8mL��_���D���27��`��u�C�7-�� Qr:�7`���p�#q�I���y��O�xem�;a='���$K
R[�c!b���c|�$Ķ6o�Wk��-�\���]o�����3ϼ��9����e-�i��9T��uK�@x5�j���Rpڤ��nWh��Q�

��:�)��t�u�� �������LJ�=�I~ 1��
�=��Zb�X[jb�;�'3 a��D���D�l2>؁WO���^�@4�G��~c
��ym��%�R̩ΪRaC_:���hpB�,�Ǔagd�9�jV"~/��6�-�R,��ߒ��}`p����dw��j,��/{�	z��+W���F�Q0y-!��;~��~�s������@*2?�B%�D\�t�γ���zC�B/��,F���l������wB�Ɲ��/5Ul�ˀ�I&V��*��D�WQ�����=�����-̅�<�a�I�ӖA�9{�Wv;bV#�m�k�)����F��]�FS^����R�����ng,4��k�w2s	=)���(�p���q�K��rO��فG�PU2��J��x�R���ܻ����"Ռ0� �3{�<�Z��G�SR�M�6�����_SUx�.Q�:��tx?m7(Cjbs4f������,�3C	s���n���PVl��+��q�����i\k~9h��۾j�h��P���7��=¶?�[�u{�R�⓿���}@tkgJ�sm4 ��
#Kw�V�^��[�X��ނ�'�x(����(Yߠ��y�=�K\=�=���MO$�2Gu7ȐPP/���*[9v	`��Ė:9��\L����.��<�OK����je��y�/`.��{e����2�Sju�K��^A~mp-� Qy�~��u`ڎ���x��ءmZf[��L.���g;�i�K����۟�k�_��Z��1���S]E����g�3�8 ��Qx�N ��
�V��ƃ�T��;@��u���)2��( ���͗==��x0L0�Ĭ�ˀe��+2^�LJ!��`�.��#c��z#�.�D����jl���q��b���Nǉy� �뭱�ŉ�Cᮩ�4�&�<7D`H�@��Jc�`�ɥd�[����]�g�3�w10�� 5�����>��GR��$Xg�wteZۣ&�%c��G�YYWD|sɥg}�*n���l&���o��� ����Q�2OI��TAϣu��Y�sd#r/��o�!yϓ%��$wgۚ�Ϸ��U�b}o:�G�'��f/=���H��;�Y9�|��y't��"y)��t�,H�bH+e����3�
u��� � }e���j����N)gy�L�5iIr2�{T��q昭�x�l3s��c�F�c)��t.�ڏ��+?�O��x��ܕd�o�<��UT�|�qs�K�FrRt�)Z� ��w!k���7�$�3"(־3��g���b�eЃ�`��'�S%�@�O*{�$�o1Q�܏���~���]9�fL�z���eZ,��5U24Y�CJ�\�6�R:'0z_����5�M���m���֞l,��TP_tD�P(�w��_�&-���H�~���)Vvh\����S93K�VXw���,ҀIe��dM��Q��Ħ-��o�����������bu,Ȭc䵅����/�#,j(�;͛�g�\tl�z�Y��	��}��~	/ic�k*L1�cL�~�Ő�q���<C�d�`����,F�<���%k��;i}�f��	�ת��ܐ�\�ߓ��>`��x]�ߥE���偄W���/�.s;�A�������,��#�|3���)�|s!�*?��!19�V���Pj�4��U�=�k�*�M),��[7=�М|Pp$�k��� �,���>5�7���@D�d�ApJ/��>h�G�88VP����M���� �P�$��EL��F��w�F@}v�w��D��6���gaG<qW����H`�Sr��r���p��-�Y͊i�	�3qb��Ee��q��������|�C���Q��}�ʌ��aZ2��� �51�3���'���UKGh��z8s4��:b�o,���E��+x�h*��o`҈�����W.YB0ˢ+�u�n�A6������N<�<�7I���.���
6��'i�X��q2��$l��}fsN�1[��{�LY�/��ཟ���HS��*K'�!�` �_��G�Wރ*���˛�S���j���X����N����0��vSXa!�fVrW��@��B#���wu9�Ź�ٷ�#vc�ۚE�G�&w�ocBڪ�apM
�0E�ǀ�¥�%��e�����S�� 9Ľ'�Zꩰ�2��%P�����fe������+̽�������q�P���P�����t�RP^����]��\}�7FșEw��S�0]h��DcE�M�ƾ��GɁ'�U*qP�67�B�.�T��P<G4�<[VE���M��dǣ��d��G9X_�lr�ۀ��`r)��3ݞ�u$�+�ll�~ʮ�Q�����lTd�T���u7��|�WY�)���MK��)8/�vjb���X����rd�q� 58m��1Y��Ao���4�`ʏ��$O�S<w����5q������ҹ�(��p��Cń�R��X��N6^�|97�%Q�C%�|P(#�q`8z�fm������6�G�r�~��Ry������.�y_U[���
;�j@�i9C��n#r����������T�sD�ʢ&�˝�����z	$(cC�4�	�9dK�J'�M@!�u8��c/���]�5�W.��^���Ж�9���?��oq�k-e�1�R��{S=��P�� zޘ^/�N�,JH�xp��Dzғ���a�[��ey�B	n�"3;=I��<��~|[��N����Cc`�u�%����U��)*5c��Po�������Hm��Y����`Z ��=`k83��*�`����>��o۳;;���Ǫ�'�+�횣$']O��F���&kk=�#��G����9���T3v�9�Gm�@�^��X)˾�a��Cgtڄ�-�����'Gvu�h٣�C�\�,������m�:_0��anf��`� ��
R1L��W90���&G/
z�RS.�րg�vj��s�0[|C[����~G`5�l�Hej٫���W@�p����â�D�~e��r��n�x_�ڑ77Y��S� C}o�(�e՟<|�Dݣ�V�9&}�=va����8����bQL��6����;�pc�tp0�.�%�- 3X�蘥��
 fWv�Ά�Z��v�u��dv@��� )˃h*�ݮ�@*��A�jXj����z�Eұ�V���K-��C�	���j�:���O�y�59�hr��7�f�F�Y��.ьt�ʝO�HT�v��L>���/`�Af"�G�SWt�J1�W�!'��B$��%C+��AOXч�$FM;�{2T�И�^�Z�<������ɯ�ȥ�$i}ԟ:��@k;�q�K��D�y�w�D��9��o�����?����6-
�ﱪ1�9Kp��h"���/i:�*�˿c�8ʥ��q|��XlxVHYEB    fa00    1950��/��p��}Q|���Вx�̣0��h��"���q�K���c�1����RS���������s-&Ut��C1���a�,S���{ҥC�b����P.�CX��ʐ򕸒�V���8�T;���ͷv������H�L	��<���GQTy#��s�QC��<��1�ǜ�Hf^F/��X��s��u���ُk^��2Z��˙��@�<k�a�aTf�
=Inl����/�Z����lVq��u���x���o�f�!7M������8"yw
�ˊΦN�%��-ѼU���D��\��i�'O��#׮BR�9�cb�%��N�4 ���QR`�]>w�{~'���5Q7B%*0X_���ͨ���=Seka�!d�z��O��٭�Y�߁y�GկOlu ����� !��㎣0�C5����j9G�+;7rcm��N�T�c�7��^�\Th+Ն�,g�+Ķ�Jα8KÞD�<��Y�yߪ���`�\�}��t�s�3J.�5�t;H;��\E�2���q��1|�5{�n�,M-\r���&��C_p��""A;�X#��XB��L��ܹp��� &^b4��t����z���Q��SOwZm��*���@��b[ٴy�>~<-j*Ek�Kn��\o	�xQFǁ��� Z�@/O�]i�5k��Z��5��տأ?��Gbx�g�hB�������JO�Ώ���#
o�s)�H5b)w��Ik�,ɜw�SG���8�௿�>�`|����ku��z�݀-�L"`�G9M�?��3�}t@��Z����r�E=��h���B|��=�D���� =)z��O�_������r�ɘ#P1v�-M�]���Cΐ��9���?Dƪ@7���F���s֏YU��z����
�~n���P$��T�G���������֎B8_#��z����%>V\�{Ng�G�}���̄-����U��e�����8,�? <�݂#�D�{w��+�{� ib�7�G�7$��x���L���FZ��t��h����+HN�9Խ�0�à�B ����Ϳ�ڡZD ��ɔ�6h!��$���� �k��MQ+-�gQ�Ļ~�)r�;Zys�ʜqp�f:�D_O�m����dz*�o:���\D�%������s���p<��.�D>w��?<�7�>~�uK��a*��[V��2*с��W�#�AԈ��ZkUY��z=��տ�����f8��W��ou$C���1���K�)`��N��b�;���K������2�D�F��tͼH�N���J��8�h%�u#�[r���"�7�Q,���l�������i�3���|������/�B�,J����	��k�}h+�|W'�<���ܝ�7��JV�8+3��϶�����/��RV��Sm�|��ԅ˨{�O��f����	��֐�l!&�%�5��8}�`�U��L�{P�C�*�:����`Flݜ��(G=QC�Zfoҥ"��â�H���8�^\��EU���PܑN�{)�������l��tV�E�?pEJ�_���J}X���v������rOŝOuP,6(Vfc���*���\�r��	ba,x(e2b�����3��U	1�Q���o���?<�|DJ��r`���C��4�n���'����7�j�韪��� 	t�̜I�����T��}�*S�^�l�CRw�!������N-e�00]�8t��6�����̚�_�� �k�u��?!��[��Y��Mn	�dp��n�
�uu�!]�Dx3ƴ1�=�]#l5�T�e��0z��ɿ����������oewJ^�������Y�<&{��@j���J�<�P�7��i�I�>La�hi��íi��k��N8����6[zw��������Y�X��
}͛���~G2��j�art Q%��1��jyGO�u ��m ��ox��R�^r;Śs�A������x�o����Kx����xpk6�}�L�w���ʈ�MϾ��������D������F�n�I([J�ݑ�Ơ�/��E$�*0�%�#�_��b�n�f$�S���3��Ktx�pJ�U'ۤL���i���t�R|'�[$*J�A�y���<��DI��R"� n�H�f"Wt�R;#�$�N�N��G�����(�};ttJe��5=o��Q�@���H;���Nc���cT��	�@�ﾎ���F����A�@@��򹛥�	�!�t8������J���oo~���p��j"}�-�D�Zw�e�9����EPf�/y[�tH���*gR��p0�>�hG,�����i�SY�9��u,��.{�6`��`�Sjq}��������P�D���!�؄8
�]
gOӁu%#8��B�A<t����"K�:�,���x/c�8<����o,�ԩ:+ܙ;A
`Ӗ��Pqq�54I�H�K4������rh!�%�<���E+���	I�oy}�_�~k���-^T�	J�5��ԯ��&4�Z���aZE�J:�%�H�c�?G�`n����?zS%���ׯ�9hLX���l>	ãH>�5)�W�0�P�7dS8& �T$�4Q)�K?��I�#SFږ�ay��i~%o}���Z<PZA*q����H�=��~����7�8��8��ƞb]eN�q�����1�zߑ�k���>�ؿd�ԑc����Y�����~9Yl�+7�>E2�@���K��;u}� �U��~d����J�l~C/	H�[(�3�����|i�^�.a�;���q��\O� 4�gH���3�����o��ѻ��h�%��޶��`�6�t�"G���}-��g)��Tf���h�@��L�t����I��G4d^]@o��	���r��+X2]d�	f���t?�ݤ ������K�b��t�m=M9��VJ�٩����s~�(�s���+t��(��@r�,7�ϥ�̢�v��1��w���Q�}����("Tz4��4 � ��� �aP�0�u�
�GQY����-�i��v+W$!o}�=Ds�&��ZhKM�7�϶�%���zT��=c�Z�o�ݭ��sV�Jo��Y#l��D��D'����/Qۭt #^ "��tHd�H:n�6R/މ��%�+�%j޴���k�v�]К���zN|�Gh$�SDf洹RqzixˍbI�b�6w���D���Ö?i��
��uu���n�sL�F�T\��h�vI�C�,��H�zM1 8I�l�)��0��p��"򑓤��!���s|�ܹƧZ� s=�T1�Qd-		k���0�9��$����FDWi"��#{If�Q��7%��N2;$���1-h���M���'~9Ć����t���Q�uV�T��>���՝F!_�N�.����@3����7�@ '��΍$����Ra���F����}I��1ZF����P#�c<�/�zP��Mr���ţ�z��ܾ��L��)>�[n:r���[$�b`�;�/O����κZ�n�����w|���0��c��<ܐ��`Bq�1�?%Vb?ٰ�_���x�q�\s�5�q�&9Y�����ڌ�xM y�q�-���򲑤�
��dW�l���u{R���{�ʻ�R���q��Ό?��Ѭ�(:�v︵�hUˏ�3,���iG�j�~Js@r'��.ׯ\�<75����64G�o���ΧnA��#%h+8�4�^�:�t'V���~�瀾�]�uN��Vm�;ȌH�}Q�}o��0��@˛�J䳝���sU������E��Y𣯑��L���y�yIp�V��B����؞��'s|j7��ӄ��&�h�U�6�b��/(�`Y����͞.�H x�&��༇�
n�D���!#w#.�/h�����c�v�j�\�|YvU�\��Ü�K.:�9<�G�N�i�]�f�A�#}�!0�h4���� 25\؎�ض&t_{��M��å��gF[2m��^�����wgN$��� �6pQ��X���o$��eZd]z?�	Bp�p� 0?i�}�AV�I��S��M��Uؤqo�((W!�X���l%n�8t�0�pS��t@�f)��}^�;�c��`����te�3�i6�W���}	�\�����nĈ;G�s�����K�mj+��+��Z&m�&�9<�cg˯��˃"�e�Y��.j`���gF��?*Hsi�_�P���t��Q�mԜ���m���U`�%z��~a��҈��D\}H��A{X1��B$����L귪�HU��?����5��XA��,��9�+���jq}�vD��XE�s���)��rF������iX;6f*}�	��#{jm4�T:|O�q<�B���r���ԃ!�JX��_>��=0X�?9-ckΊ�Ԅ��9)	�j/?�"���H$����pH�<D�Q��6vs���΀���2ڊ��l��e�Q�ܚ��8)f 5bO"��Ub������9O�ۙe��ʫ��/>�׷��TD�,���5NF=�0Cr�F7�#o-4�4�/�8Q�g�L���x�����½&����� OzT(q����nI?k��4B����|��Ixq���u֧�O7@��6�*.wc>��9_f��������=�`���8�V���2r����\r��F.�.��`Y�k�Z�?���=�*�]��t))m �,>�X�V��G�=��G0ER��G�ǰD�����oG֐���B��D.$x ��3?�^Ǟ/`�2�ʕO�7Ї:O67�TS���p�����6��q�A���K�h�#�|�v�T�+��k��V�؁�(��J�}i\�P���/�G���@t�.��OT�W�+��"��n"C�(�W�Ԭ�,�3�Q��5!A�-@L����@��F�ͦ�v��k9�b�B$�:�H�֋ُ6�$~����Fό�J�pL�G/��-	g� h�r�J�;�X�< ���Rv`+NPC��Yz�����f.����`�5��<t�ן��{rV%
E��/�}{)}õD��'�+",�z�����m�i�;���7`X��|=���V%Z�;S�|���	�VA�p~+KkK��|��"�ّ)�[�ʁ�8ʍ������kzs�	�G�ve��+tf�����pO����	c�@��{<&2��Vʧ����y�P�v�=���d����p�%P�Ι�Q�1W�[��Mu���7Ol��9��<x�8� cZ��]O焄i��*�E{��p�(i��F-}���J@'<(�n,���DK����J�{Q�#����c^Ph��;���Wé�W��m�-�;��+i�^�F<L=�Td4x���gRO����R�a���F&�$����yԯc|�Z�&����N�\(�E.h�#w�8^�X��%�����ꁐVFO�CZ��۽����W�ژ��g����FU5�df���0�f�Ç�}_I�"ݘ[���5��<C6N:���*��������v-`¡GK�z \��Q��p�k��ޔKm�8N}yd��dsmem��-R�u2��z�l�.��IM�gD{��x
D�_�K��t�J��ݮ��Ɉ?��>���<��富/�=�Q��>ef��o#��쁪q�� ���V�{yY��K�i*�LiuD}�H\~F�R^)ഀĶp|U���TO��Z���:8���;�l�C;Ȣ�U9�t/��x�v�Y�2��é���a�-��_�q3�,��3��	�V��|�������0�y�����8��W�ܝ<+
#�C���59��q�vU�ϊ"2i���y,2b��Mˤ?'��#��]Sl�t�J&M1��4�f�i���;�+��h]�_u�r�:���xt|�T:��f^��,����,@N+�X�|"�Fa�aG)n�įu�a,����)dT�/4`�s�פMT�SF��+�l��:C̅PG6tda����BF?�__ڵ�\@�11���7�1����GT�Y��T�D�s]�c��t�?fiFƜ�s!9�j�C�9T;�8B���g
��L�KD��:�t�e�1<p�߳Wb�j�æ�����I�-�n�B��c|)���o����E����qq9��B�����M%l�ϯ���˚���Y�ih�kxi�����Z���³�P�$q ��0��n�1���h-�͏�J�{E�j���>�_�����X<� ,Ň�
��(�7e��O�8�Q�y��K:�vC��L�[߸�f�	�nA��q��-��uMȈNq<��܄쒷�W����f������U�:���p���d5o3�d(}�؂��8Eۈ�P(oy�l�)�Q
���(25��@1����n/m���?��c:����n;>�i/8�[d9<YA�`3�b/�<�NH}��|�&e��$кԼE��X�LH%.��ΚW�XlxVHYEB    4f27     d40����nm�$M�t���]�!}�0��=��z$a A�QaŐ^Ћ�M�ޣT�o������̠���K/[�^�F��epF͆|*N��6�*;S٧I�=������[�YTAY��:�t���t�Fg<�[d!��6>q�u�Q3�p<����Sq���	Ym\	@�5����#R+�e���ҍ������&��	U9������<��m��Jl;G!ɷ�
-�ASw�W�*a��7����+7� �8� ���:�D@��4B���3�'���F�u����C��,�#2@������W�����#��4:�U(��
_Y���,)�xi����p��sw�5�u�̓�ͱqS^��Q[��bĐm�x���c��uSh6�f n��p'��:S 
C���?n�ң׮�G���[�\�X���J�m��7ŵK�aנ��T�$��P����gf��n?80�c�҄~~r���3�h���~���k�Z�FD�G�e�x^E���q+ �Է�4V zˢ�I>]��$�����
��Y��� �Gة�}����|��B���'�������b�?�q%�;j��Y+U�w��,G>t}b u���A5�PsĊ�Ϭ�u����'�����C�|���=���_�hr%�,�l&+��^��C���d��[۹{8�s,�Pd����E�@���F��`K0:�ݵ��0�O�H
0!��2��O:/���c/���G�[�JI��SK{>���#���z���l�k��y#��P
}}�ݱ�6��+jV[�"нI\�cZ�#�vy��y�w�BYc��_����mPE{�5�˒:#�q*Lտ��=�vۧ�C���g�P���j�򹈔j-6�W�7���K�F���!N�\�uL_f'�s�C~<)�H�u]��wy^
;�A3(o�5k�n܏S��lx�t�I�zT��B�nJ밌D��;:X�w`l	a�����\B����>77%;�|�#D��D(�lr��py��N��u��\|��+U���Sz)�#��CKB���-�z���������^�$����ݺ�Ὲ�)З���@o	gJn{7Pv�:9mw���Q����̼���{�O-g^�0i$�ʠ�&}�[
�c�Jp��S��sI���>Ǣ���V_�c����Ch9;�Op���x}ś8�d�L���V����BXK��$��a�)�&RV\�3��M��}��zȨz4 �"�Ӌf|�����iZ��ݚ4���O$�����ZV5�������m��Ɩ��ѪK�f�A+���m#5Z�r� i�ƱK�?�zl�k9�k2�܊L��V�c����3�ռe.��o��9�d��u�����,Y��x0C���x5�ol�썌�+�l�9�p��#�R�;U <K��03ˎ^����_���2�D�t0K����ը��4���:��w��W���*�D��#��P��f&��U�q����䶛S���#ǈ���zXvQ������l�`��ƬT�d��1r�¬1����T��Xy��sZ��	*�㭞b���+�^-�Y��ʤ�0�h!tU�Ņ ������,v������Sh��]"��q�a�E P�9�$���|u9��J5����Q��Iv��+�>��s��0<W�Gُ;6I��.=��R7𪮍��e�␹���ČZ�.4�["N��c�!�D�q51Uk�(�^�#aFj�ƳO#�f����UB��콴��顳�L���$�,]���N�
eE�ƂE�}����8���:�b��i�M�49a�g�$c#)1v}���=&E������P���/LZ�����ؐ��)�\�k`;1B�B��R_/��'�fk�v`=�t�?�b9N2��	ByJ���yĺ0�%ƺ���~N�<�� ���8�y�ǎ�Gҥ�E �5�!pV�����W��"�9L3.I�ؿ�Xũ����������ި�:�E���t��@Q��An��<�uS^ kĹ=�9!�&�W�<fc�ґd�!.��e�Z�Y�^�a�c���H�����yn��uz?��FU�� *�(��OY�m#��[�ә��Z���al��w��-�\O�� �%�b���߽����~5/"^�Mթ�g�\�B��F��L:2��=��zB20����/�}p�b$�\�ZL������Z�ߔ�騈Hj�U4)蓽�� ��O6�ɺC�c�"+��GO��*���.�X䷰d�H�"��K�>�gHf,8�$;�
fo����ܠ)"�.Ć��k�+�7��Dx(��	A�1;���#����s�EϹ�PQSԤ"�Z;(�	jO�R�`�L~C��&f-݂�
< ��nA�^�\[Pjl�����H �\)�&�!������^�}����%@@�[�ahts�kupv\!bA,b,葆�+P��-�N%���Jx��q�����Ճ�]Z�;����GE�AGu&���Lke�N��l��@��ԑ��j΃��z=(Rl���Y9��P�@��f�I�)6"���}j`�<���d4�9A����&y�r�����4��G�_{���p��A���Q/�o1��1k$EN��'��x�z���
��S��P�˅L#>@ja�`^Q$ �SY��������Uت��HC�qZX0W"���Oк!��z-�B<�]���{�}�5�����
-	�c�nQ��{E�с�,�à�nQ�g��DU���8{d�m��o�����ݱ ���Xl� �q�]��F�"D�je� ��.҈E\;���a'���Kݹ>��(�Q��G��˼��+!�w���;ڑ�s��KåQ���O��Vˣ9MUX�A�$����G�K��$��!`5��Ԛ�ϴ}f=���tQJ%���2]?#�\v�88�tB�
]+_�X��^�$2A|<q�A���w�s �R�T�H��犂�24��*�x�B��v�
��n���}ٖ�=��fR��j)�'a� K������P����Ϗz�Ǣ%$'�L���&��~�߇l�c��|-����Ə+�GY��h�2�Q���+..Z��<W������o囷�0Q͙�_�G,��ǰ���,�1���t��B���J���4����^ �	u�'�C�F�I>Y�?*&+ ��U=��7;�"RG��N�������2��UUP�əd/W���X���}�d�F�rD������k{�>G%��\%(���	��if-7�9�f�֎!}��d��e, x��6[!�ׁ���T�(�l��R��h(^�����CYg%ػVt�Yz�z�0��f�,���H�A��~؋c������9p��Ұj�>9�