XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������J�=i%�pC��s#�f��6����m�TYǌ���sξ{7g��}�~�lb�ذ���K]��Wn��W d�0ik.H�N�c�!6�"W ��]����QQ#�Yz�cP���5T���)%�뉏]ihv�Iz����R��l���Gg0]k�3�uR�+L�T���p�@���5�&�A���5�k�#�Ǳ�����,^,B]߁����������X���z��p���K�������=]��c(�\��T=A��B�L�����!������+�!o����7R,�U�l���%�E��
XF*#�8�>���!�%M[O��^���i(4x�lԫ�䲤�1+�>�����@C���<D�0;O���@.�� ���9X�n$D-���hl0��s���M>�ќ&ҷq��c��a�h4�-�-���,GF�,�{�å��uad�lNx�N%sf&SLḞe����@U�3�}"���2j���X�N˺m�V�|1��w� �H��E�f�+��:\b�%N��lݘ�k�N˩uc0Bf���}��axB�#߿�Pd���U-]�J��EId�X[�\B`X�Q1���D�K[s�G�*�	N�7��4qaICl�X���<7ra���2K�C�� �彃���H.N&(f�	�*���������/R�쥺|�uj����G6�6<[�d1�l�J��٘�ѐsRo1���+
v���,C�S�+�����U�_�W�8n� �n�16B�,�y�2ﵘ������HXlxVHYEB    3504     cb0j�y�j�)�&O�#ǔ��2�('�{�$���30=y�Fc�>�I2L}$���Pm
���c��2�]��i��'�������C�se�;45c[-���w��Z���k�M��ы�=a�h�bn������tIv�����qGiT�"�U�k����5���hZ� �@�l����dɛ��gdO�]�4�%�6�|F'p����~�&�ghpiÊ��d��\�,�P�y���9�`��8������&@P�w��/�_��o?��}3 Ɛ�lX ��`�pn�]�2��9�ڇ�@e�)��,��q��=+g�B����ղo?��1.T����y�v�lz@�Q-���L��Oϭ��v�&�>ε���z�s	{�m��Cgn;��h6��I��F3�����)��p�s��lV.�b>�B�hFd�s0�֘Lo�h�P9v �Ʊ�#�7���}�x�l5{��9�Wl+.�ʏ���k���q��o�i3ԗ�1�QC����d1����u
��� �ٸ���x��mT�Ў
�?�-�A.e�*�=HР�r�AZTUV�͋,���R�Pw������3�y�A�����%Wj���&��0�O�ɣX�պO��RoI����E[�^C\�� �lT/�;�>����E�ňl\�f9I�NG���xH�AF,���]�z_ R@\�R�]b�Uz�T�~���og��,�9E�vD�h8�,$�~��28��7�s�:�cL�˧��g$�����%���\
�D�����V�������;h��P�t�\�V�z�!�9(@�J�Jhf�U8�������+�%�xN������yj�	���x�\p��0ShRnR���0QZ�`v�^���,Wt��&�	SB��Lv<&S��Q�HAD��^jV1T��	}���9��E����f��溥�>.z�`U���Fo�IW�ѝ�O�%����;�3;F�}��/�n�����.�����ɣ�U!�T����03_���{��+}R�t��(Ɔ"B����Qv[X��V*9s���U�-n��.���<
���Q�� z"��#YAT����$ÁQ�O����hFS ����Ǌ�T�Q��o�(*pƐJ)An��Sr޺L��D���ʛs`���\����2�a������▌�z|ۿ��c�^�����;��B:��������L9��!�ۻ�dJ��e�[n��Tc�G5�sp�����m�t
�yU]�f�,%�������⚘נk+����芻j��n�j�(cn�%�g٬�C��D�Ł�fq		����1��Srr�xK;|��j�n9��2cBsiA'㏻�%�iX���Pan/�d�ݾ�����<����גR%M�.r ���!�S��Z_�dvi�X�LD�,3�W������`���h��v�����k�g��Ob�d�l;].��#��	�"�<�[ײ��\
(�PʦmnĒ�Z��Xf��D���U;5�,$͝so�~�5GO3jYioBٞY=&Y?@���5��d���
��'GU��Y��O�p~�_��I���$;���4V�$��c%	���M�͢�Z6)����$>|�ސd��aNgh�	�\\m��E��*�CM���K���ӯ���J���Yg?��!�}WلQ����nl��� �Z����+��R��MۇV󮣵�1��a~%�f��V� �߲�S^���+&��6��Gd:�g%�Ev)�I�M�k����k��.�1�S-����	�����D�%��b�͆�JL��
DѐS{�z�'���ZA�(��\m� �Xc����G��k~|����Gk�Y{����`J��i$��@āL��r��f��RU��x�T�q�(]��n-Qªn[tE�ʍ���ӵqdѱ|����J1��'�9��]�a��6�M��η����:�f��d���Q5W��q����Ύ�8H{��?lyՉ���#�7��g���P�hy ��T[���Q�+��Xs 0�ԉ�ي�B���Y<b��jBC0�3��Uf'w�W���Q����2����i�N�h
?7����p�;^хmwT�ƪ�̓��U[�\�V����v1n&�l0=�%�-K�����@�|��S�Q�\|�c�&�J/W�cP=����Y�uיm�f�9���>�%5m�N���8�VJ�6u�P�F��+��4�ugN-�1\}z�'��KE r��BG�0�yH|�]u����
�
b<�^���CRl4�0�moT.�I�YSҵ�}�G��=)�[;���u�X~��2���u:�x�'�D^��` )�km)-�����, h_eY��>��a��u�䨿���-�wщ�K�4�Ur�B �͑�5b"��̑��B��)�1��a��n��z��5��L�ϡ��ipl&&�!�ܮ0�o?Y2���W�ih'GG��*�"k�}�2cOeWP%��*_��W����Ů�m�X�ϖ%����Of[���{&C�B���O��[-�d��s����$%�_��o��s�:�q�����ת�����HF���o�f)�1�;zJ�5�*���!�ʲ�����<��G����Q#�������q����ݎP�)�ȫXh�^p�jg���J���/FY�f�����;�q�����bP8s���y��&��`0C�vȁFcg��竛.;�*�^r��@n��#�mq�˩�X����=P������}.D�f��^�)A�λ)������D`���#Q^��͘����kb����(U�}�-R�V����Z��T%���!�F�9�j3w���$]�54���Oj���y��G�T���Rj�H�j\S����}V����_�:F�ȶ��,�g�,���>��5�6H3Ǩh�݂�	�@�W�0�w;�Y��eE	ި�t9��Ѱ���<UB�:����l�T%�53j�ar)����9�����3Ę5���tv9ұ�L��v1jKi�"�I-��t��r\Z+��6�x�}c�H;�8cmu�	�>޾8$ޑ�GAUQ�Dp�G��34Z,�z����VH+ep�K�����蹫���� ��PEc�����9��4 ���*50d�[̅ +�[~b�ȕ�3s�K��"G���~H�߯WwČ�zT�x�e�1.=��x?��A��Ez$�c� �21�?�3˱�~�|��eTv���oE�>��uۏA/�k��