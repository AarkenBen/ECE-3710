XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H��s<%/6Q���������n@�QO&�I�~����g���4X�E`G������Od�����,2TmY4-�,n/{��.6$���<�n�9�.����g}p��:o#L��;꧎P>��̸��%�$��5\�T�m�:;����n�Pة�����1�糖܃�u�� v�����;1[T�ӎ�J	&F�DE[�l�f�zhVM��wO�V��	8�Ws:D�	#&MO�ʶ��%s�ل�j3���k���-����q�L�_������O��S �e��)�Pm��oH��v��թ8�!3�@j�?];�]!�:�׸%d���W�|�GKV�H	+3��C?:���_^^ �������T{� < ]�e�}ٍ�.u���=Ҩo���uz����{
�VHx��u�\�s�i��;_q�Z����3"���R�w�|ܖת&{(fߐ�a��I+��%�$������YU� �R�U�kN��"��܈�y�ƨ�H/=M�K�Aڧ��VPI8	K(�l�!��[^�\�Q/wzR8t�AP�X�`����Y�q� �,��F��r�A=�Ie8��O���k�o�!��E)X~�3�޾ߑ��?Ʈ���Q�+�mR�L-�θ���4#��CbhӖ#W�þkBu�G�g���"'�A�T����W���zxFDǓǚqw��H�>�#��	��7���-�2�����Codq�֩�����&h��J�.'B��k�O0������wXlxVHYEB    33bd     c90�F�I�+���sh�����'^t�t�3y~�������v�=z�O�)�X��M�]���G9s�o�i���}F!�����u��G)�j��Q�o�+��%b�3{�ni2�U����B��:��ҩ���H�Id�^ ���@�[_, �=�>�JU��S�դ���KeZ�����ӎ����~�'#0��;y���e�d*FV��;�ҳ7��!��y* `a�dWְ54=#��5�3<���`b��c7��E
����-9�]�08�57ݵE/�P؇!�O�m-��X����U*���C�0���q$�F)�:�u'v���G�ӻv2M�S@�v�`T�1��.����ɢ3ʽ�%_���;��	[���~�V�{!ɼ��7���`O��Z�)�6�z2l���_����ǖ��6�~Ob�3DtE�Eg������'o�eQ���.W�H�F�
� %BY�t���2����ɹ����	w;w�	*}����l�|�2�3 ����˱���G�En@;�
���f��v|�
v����s��� �~�yQ9��@_X��]�+CjZϳ�xb��</Gd�Qp�sQ	G�A��հi��k���\�����L�
�"ˢY�T��]�rz��ľAĤΨ��㛦�3��M# N{R�\2�^̴#��a6���oʺ>pX?�Y�7?_�5�����:R���f��v��]�Y�0;���j������u��ѵZD'ܹ��,�4��s�Iw�������&;�� ���'2p~7[��XI�=�i'��@�T�ST<�981W1���x�o�2�^n�E���c����Ji�Ъ%��?�J�I�#���Bq�o,�p�\�{x!�t�%��|��͜,�N�
rx˦�i�k�"4A�f�%���zi��$ؘ�iS�D�8j{���B�we#��&<�h�q�����A��#stʧ���n����+�%Ǉ{$΋�U�H���L �7Vax�df-���󚳙��[Ӷv����z�.(gӉ���9i��LH�vɅ���T쵫|��K������`�FWk'��")�8��WiOl/Itl�ob�L��مyK�\p��w���H�UD����4J ��� ��;l������7E��gu/d�n�J���c)� �߈��A���{ȍV��^�B�A��4zD2z��g��H���ekt�QJǂ`�.H�d��%��.���������cr�t�6u�b��zm�@>����{��I6����ԃk���ƫx��]2��HX	�ݩ�3?�(�Zl+B��:��+]�!Z�b�����=�����_瓰�-���$��~TLʐ��^��Q����w��m��یf�����'���#�X���$O�r�kv�6��]ߖ�$�f��;}���e�?�V_�+�>?[��k0@������#����	��d$b��-�礙��Hm�"6x�4�5NOh1,�S��lG��ƏbB���CZ'�Be/�VM�E�C0tF�n+Hr��r��P�U	{[9<�]��#0�4��E3���Zc�Y�BT�.�5��M� o%��">%��N#�q�L��ȗn����ճ�����&)�C��̛�6j�wR,R��$�r�/}�M���0U?�煷��3�G�x�^V7��������F��;h�eA�p�{h�U���>�R:f/���q��<��{��o� ��2o+��n����t.R��m�样v17�'�a>�@�W7iN�LP�<�X[�>���v���x��i{:�e�a �N�͎�{F�����x�B�L
�d��Xs|Ki11g8�>�AN���X<힩�N�G�bY���=U�#3�n�&���9	T�z.���_�i����*���˖����[���qdS����ԑ~&%��m)�ŏnD19�&Q98���ˤ�|�������wC:l�h$�
�$7���F:�΃VXjj�2>�e�����c%Kֻ�Wh0p���6
�=	%�d?u�E�C��i󸞋aEPH�}w8���*&j�uL�Kb�M(����-��F况�!K�ym�Lٺ�V��m��(��t��?����i�(�gplz2c˄)\b�����;3�,�>���e����H,���-�=J���(>�K�٭��A��J��i�P�5*�����1��S��T0��v���9�z9K�t5��cT�ܑ�'u��I�;jO�D�E���%G`ͨ5��vM���N�]���� =䓟On���s�l�d�cq�ݨxR��{th����~A�ƹ���r�d[f_w���-�ɘ���ٛu�q�����t+y�Ђ�ɚYI�Ź�p�FCp��4f�Kc�0e�Y'L��3�b���6���6z��� �Z�������/�7q�|Ǩ���*���<�x���͐��V�[�묙hT2�p��J^�;��6 [�X�޹�6z�("z{ܚ��Z��M\b�G���Mv\�:�"�8�F�Zن�E3�y;�l\5a�rku%��Ç) ��U��F��Z����)��uV�Z��Е��Z��r�?"��Xkrq��;p��<��M{���<�S~��,�APg��]sK��-�w������Gi��������	`���,N'�5A��횧I�icR�[c�Aj�m����F�,S�ۋ��gbO�ڸC�,�ko> �W��0P� vZl^鰪����Lj��:������YB�z�9�:�`��ijB�пO��eB7�ք9K)�N�˚	S}���D�󓟺��ߣ�=n��0YU`��W0t{a��.�+�R�[�W�̼����}6�;��h��ٲ��7���")���*>_�@d�'V;�0�B�����H�7=]���j��*3��%��}�]Q�@��61�,*��� �w[ɊH���2c$�(���(�q́�[k��\5ۮ� �J�1�K��5���B��9�G��-���E��jgRmjB�P��4ǡ���"�E�d��Io��\g�^J�ޓR�ϣz����"6�	%�A���&L��I\y.2+�������	U*@����q�L��!��nH�&!�,C� p����WaT�H�A?a�S���W���Q��!�+%�P��0�u�k�·���p�f�s��M`�`f���г8^�w-t,���?l7�R���