XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F*�e6{Y;[����ї.��1�vz�����x��鋽7!�u�Z�|�OJ������m}^�D}Rl��^W��zU_���Qcl7��I���n	8��m�"�U�)�i���NXp��^�_+�Xՠ9{��Q${����3W"v 5h�oO٩�w�gI1>��G����N�idh	�%1W�9t�e$+�<s�����0�B��T�#+����`�����U���Yt�^@���}
(:ќ4�\NG�}x�7������/4�%��UX��ϑ8��%�p�����q�5`CB��,��
�P0�,M�T�oi�~2]$��5�,�*^PP��h������Z�:�͹��e�u�=�5��������;��Ƿ�����^�̒���E�1pU}M���A�mG��OS1;;]u���/Ɲ� F/ZX>q���4�l��BE3@P���)f�)HR���N��`��� Է(ϟ����0=o�2o�Ԥ���i�Gv1w��.�k��ߗ�?�-�ⱡ��ڵuD��+k��+�/�Կ�K(�]�.�33�VK>r�DV:w�X���7� �s��qZ[�M��}$l+&H{
 ����t��|��"DD
��˟����o�G!>eyC9<� M�/�V+M'�%j}�l�{�T��+�P蠾��J~O�����h"�Ɓ���_Ƌ�p�6���i�j�x�r�aQo*�mG�bA7����4{�_�{,9N��(���A��H$��ě��1{�����7JD�A�ɤgXlxVHYEB    9efe    1be0����N��u�\J�C������#���?+��En`%6���}oU�Yo!���aQ/�d��+�l3l5��//�ii�.�k����������ʵx��<"��2X&��Ѩ��)&�9�S��g��5��E�	�ӝ������9���A��*�	�������e���|�Etz�t1����k� ����n�s��^�3� yD;^o�'��;gTЩg������-����:
�Pk���Ⱥ�������(�P�fҝy
�{;L�A�߷�����޴I+�6ޗaANS6��mk��Z�o�h֛���	f Rؘ�J�j*���e�!����c�Qe���0k��kC{~�s
߅
eIy��:��x�o]� ~+U�_u���@��Y{�>�*x�4�Páu�~�p��mwwfV��0�9���&О�w.&�@��9��� \c��!���Qmn ,>��F� 	�V�����&�r�I�pv�9�S���߅���3�6e��fK�ҽ���;0~|'C��5�$�
P���f�RY���blr����Rq�m6Iva�O�<����/Wy��M���^�m��äjv�8�-]w��Y�-��T,7�/�	�Fk����m�Aca$�= >��Ŭ���(��
�/���T��Q|��٣�?�[s����[=A��L���*q��ݿ��fcA6-�7<�#�KA�;��s�9C�aץ����X ���k}����8VD��p|*������V�n��(7j��A�p݃q�@�I�d0�T㤬�C(J�H�S�}�(v�t��P1�_�H���}�
����.8��.��(�s����|��R
i��g1u8ɹ�i��IX���T{��u2E��MHqH�B;	W�� 6S�̢��3�0J����퀔X㧫kϱh)����8�ʊY��m���tL=L�R?D�w	d�K2D��P�c�t�D������J��ɣ�B������D _��y��!#��A��v�}���#�6�����`8��VTk��R8r�N�z�h���_��a1�=
"��R	*�|��}�f:�����#��:A��8�3��ڊF;m��Po�.d	�,�OS��~k%m}T���Ҍ�Ct�XeP��[�*h
$ý8�6`�i�y!�$x�4�x��0W�J��[UΟ��cP�D�漗.tn�Q�!�Ƽ%�$
x��(��",���-�(΅����!-�|�L��I�M�\!�,� �I=�x�K ��V���3���U��a�+�i ���c~1?��Zƕ��S.���B#��I��Ms��F�f2��z�T�(��IȻM��6�|9���㴼ݪr/ ��"��z�l�����U�)�����=E��>��!C���{S����<�Α�}��/g�Q�&(��W�p�_�P۶4�+f+����[��FS�֮�h&�
4��	S�����-��X���ބ��l�M�����>�I�ɦԹ����A��0ٿ��{N�B)��H���	�SL�jT �(UpV�/	{\W����5�h�x���6n�.I�!���S�&�pǿ���Z��"j��mэ�Ӭ`b�F2: Brs�D�[�b�mK,��Tg$�+Z*0�0���	1�z�9���x�M���Z�����)�������p#IE,�Yq�A��ALftu�)!�4a����߸}pk�B4���B���w��K��$��jTK�!iUQ�ey�Mס��� �[�!��.�d��'�>��a
ƚ?�شp�{�A5;�?�i�4�W�e��L�2=[��L�T���ƣ�X�8��o�ö��.�J�sk�R��+�H�{YFOǼ+��=�b��m�<N�;ՂO�\��A��T�A�ы����ftW̪x���.�����z�[+\���Y6_��D%Ѐ�f�8��m-X��j ��u�g����mg
9by� p�k� �B��Fɥi䢐�B����~��K�	�P�:s�)��r�����/Y:N6lZ(���e��ID�E�Ȧzg7�qk�'������'!C��|�+��-����
x�	LSFS��{�o�\N.W�q$�џVI1}16�#Y��IhϬD�L�3l���]��t\��3tq��2�j�q�n�q*��i�agXԩ��q�����C Bn24�݇F5����i��U� �T�u)Č���k~�\�Δ�ڙ����닺�_y5����ٛG[��=��a��ʩ��ɭ\��s�
#�0�P�W6Zc,�ǖ"%������]@b��}
��d�,e�/x ��+k��폃JE�\y�4ԧ����9|#Aɟ��Q����LUW�GW�ПOd��y1�\���u��΂#�H�#.sB�D���rB �o���Yĝm��a��#��*��k�K��#������&�pX��l�z3�ؠt����ҟj�n�ؘ�y(��UM6��c�<�DH
�C���U���Z�*�S��@Sҝ����Qjp��\Ug966�ǎY����K%t�?�M].��n���g��A@Բ�É��u���<]���U?���� H6���)���U�ZC^)_�	mI> �8�5B����*����_����_V�;�� �v�G1�3�H�����1�Cs�.��m=�K��zh�lh�E�ߌf�J����uD����FhKm��YZ�����R!��"�Yu���	X5��Fܺg*�eI5k��]�O�K斡ܬ?"X��o+;4����M�Sd�^<��}��+���k����6��=n~�N��0j��jhx?n�#�եx���Q�?L�b�0��7���R���n`�lC�|~�{VecMP��t���&Oi>*�������� �Y���ķE �`�����S���Ip{��g�/ea��{��D�)��l��7��3ll��k\e ȓ�C3]�~�C�.'��Y�$JTVƣ�yӎ�"�caeсi��
X>�~d�^�ԁ�h��ϟ
4���]2
X]KśF+Yt��Z��?��"ߎYR�>�uyWH#���_R�3&pl@,����`���`�T9�|ֻ�5���pN��E��`�����c�V=p�J�m�������X����w��Ϝܞ�UAU��c�pd^�)�I�E��=��u���ѱ�?�O5"9��f���9���KD%Z��n��]z	B�&-�Y�dS5kNv{��á��\sg-�+׏�e�ކ��MS��f����Z��k�o�1Q���N@y
�U�ع;�6�-�7+�������y��UP�J!��h�<��x1���ji��f�t'|�{��FF� '�.����[4m3�"|���pE��Cx��1`��AQ�kF��FtKܺ�|ʘ?�1����O2 UEQ�e�6�F�Qo�jn��c����]U�X���/�{y#�)�*�c��o>��w���G���b0d<H���G��Oq��U
K]�nYef)�n\<Y�4O8�x��c�S	㭋�#O��h����.�ԟ�$��Y�㼀G�3͉"Ҫj�׺b�k�2�ir@��Gܗ/�sĴ�Àh|�,�Z��Ő2��D�"��btPa��_��.��9}+���h�uwv����`F�Xl�`���Yz-`���o��[^n�IqAojyh��`���3�[�QhcХg�m'dǟ3�9!�d>�v��@p=�B��)7M|2ꙧn�K{�A ����krk��|����l���<���7s���~)ct���<��T����/o�=�\�_Mh��v	Nѹ���jO0�S��0���q��'����UB��l&E͐}�ƌ3�!�_k�	|��ӘC����܅>��m��C���ɵ�N0
�J���k�oy���!��O�j�!�`�>���>�^B���ƫ��?�)�XC�V��is9w[�%�-"w�$1���k�j��/�@�5<xOr��ڌh[8\]$˖��\в���V��-���9��k���M䍥况6�~���oꮽ��A��)֧�P+����jb���jE�i� �i�F� �Z0/�A���BGۊ����������E��=�R�m�-���~q�B�QcB-ބbo�&��|���C���)�`B��֑=��|Q��'nd!!���8�Z>^�պu^�C�(�-,7S�WI��َ��-r��84�}O��)t��mk~���QŰ�F�5�8�u�f�����D*j<�e��v��vk�{��=�,�rJ�*��U������<ä��|I!3�5C�Ӆ�C�r)�%�W��t�ɬ�r���6	�{�sON�����Q���j-z�v[��Е��HD���Jɘ��U�b&x��c��7���9�����	�%�8��b�=7��p����WG k�C��@��m��K���uL�5��f�"��6��\��Z2p�PI���y��T�j�o(-��Ӆ��6t��z�dbHX�q��x�w��@ವ�VNְ_v4�i��6������G%��e<	.j�DѨ;fm�K�줫�,q|����uD��p�n�@���]^�.ֽ��p�
���9;�-�ٚ�*i�(ޖt0��oԩ��@y6�1%�o]�_�;V-=bL�'���G�@]����^��h`��y`׸��8;��Í]?�Cl�
��)��6���Җh����\�[�[S^��7�HXRzXhe����<g��k�[|����CV�(���y�]�TXf��������"r)O�F�y���nS:�=�ڼh���V�\��>C˗@��V��/E=�Qf1k�s�^��>��7�&��r��8o� �1_3ùN<���F?I,�-$�C�����J���`3@�OZTL1d�U�`�"U��/�hI�ϗK�r�_T��.���ޒ=Mb~�uO��W]�>������'��C��~A&׻���6��_d��yge�fj���u�L�a���>9F@�pwy��7G��1��Z��2�*	��-(��k쏟J�͜���W�]ϼ�PԂ7��������Z\�K��ʷ2����C�X/[7E'$��nU�׮�v�*-FN���UX۠F{l4�[Z��1�����Ž�,�X��-��n���jw�4�!-��AM��4;��Yvt�St�ܶ��(��_�$n��%��v�"]$���v�j�uzyqG`|�*�2���=b���P����Z�V�z��6��<{cb�.�Y�:���{S,[>��L��_1{Ր�w�U�i�����u��`�iZ%M����n�k&:0>%^��J�8�Ͳ�~r����=e��L�g�iˠN\�Vb�*(����/��*x=_RPH*���k��e"�3��{L�Q�_����?�.���6LL��f�~	�:K��s���܂h�IIw�i���Bt�'�������!x�qΟXB�$쇐@|E]o� ���t?T�}��.-�{w�{��<w��8��2<��B|4�7E���5UH˝�g#g��94�t
�o�"�p��(���U�2�\WW�� �����b����@E 
h�sq���[�3d��
*��~D����r�f�dL��J����AWo�?l�/�zIԅG�$d*U��/n$��j�ȧ���N��Kw\A�=XJӹx�ժ����	�XRUD�=�|��HKw� ��+@�F6�{��(�_A"�]]@t���������p����6a�/qN�-�׶�(t��N}h�0c��8���S��-X�8�Z��ᶅ9��Я4����
��;��374&ZX��s�{�r�koj��޳m���۹΢F9q �x�|g�����+�U`��������Yj'���-�.'���B�|��A��v�OZ4D:�����}�Ȼ�����p��"K��߆s���CK���B�k>t�I"\�á��H]���J���4J�ɗ+�w���-���]L�|,���l�SA�rm�g:ܕ)xNp v����������ЌE=���!�ɝ�x�.��B_�!�SȎ(��@~�1��H�o�%�PC��OH/�e�0�ak������E���/�T�R��#`�~�ڼi��U)�xk�'��8�@n�	��w��@������:4Q	w���q�$ca5 	F2�}i���&��?H���A��Q�fֻ�����c���j\Lf ��Z����q�g=�����/�Z���e��`%$�;�����_�2l�{O���k��t[�E?���^��ܴ��֗I��1�x`��qa�z���^w�ź�:���.�����>�ݧЁ���Wq�w��x���R�P�'���E��*�Ui<��r��E��|Y��d��C�� �/���J�A��H��� �bU/���韋}U�ZVu���)��k�"X��2����?5w�:��0�Q�H��a0�#�b�h��,R�%�j�4��K�����Ę��Z!z�!�`��-��`�ͳ�Ug�lן;n�ѡ�����P��Tz�Av���s1��5hהm`��ϯA�(�9����mٟH��뻞�C2i�8�kWF+ȕ�D�ߴQ���0�5:��|�r�pp5�8��r�PE1��NmQMv�י�|C�d!���&��6Ӑ�V��N�Zr8�o�������k��pgn����"�Js�{��{ɂ7��j�ץ7�sh-A/`�S�}�\�k-��ߘXIFщ7�����&.Gͅ����3ḚlR{��Zt�����ۛ�� #�ޅ�Si����F�(��e��N�ˏ�mcL���DU�ɨ�`t1��]T*�l�����y7�)���y+�/2)\��S��Rz��k[E���%J��bR\�k���]�@��CU���[k�?¼ا`�u�v����8<}R��m'��J�ۊ*����j��%���U�_�]�U}��u�@�W,x�Wլ�����-M��L j#i?BU�h<�A�D�g��Yi��$��4V�3J�׷�#���3 կ�a?��#8�U/�`t�_�L��EU@X��*���Jw���Tڀ��:ءZ�Y���R��j'$�>�& LM�"�g��b����+M�X:������Y� �rd�cY9Z����\�x���x=�D���