XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7�a��ia�\��gp{��HܥK�n��\L�Ɲ�̖E"�ִ����y���g�D������;	��*t���z+= ��i�￶�=�n���*���F�w�}x�
�'e=�E��T&�
��=�X�I���o���[DY�c��X��u_`���ξ��D:6��9�	)���՞�Z�v��<���8��Bf���z����F� Ou*��%F�4*ܯB�\j��["*IC����φ�����d����}%s�h.�J�h�|���}�2#
I�Guܰ�-��	`�j��KFiu2*�l�Q8�!K64����� �r��_���$��b��ځݪhu[x��"�3��j1Y��`�2L�d�Ө��C0~Є ���b��!�R�H�MR���8~�w�4e)��x�j�	�8+����>��tH�b��l�\��!\���2�_�����L!�l3�������#�y�`���@��R/H�,�ݚ��%]߅��ИB��w��Α��/Z��PqT� ��wQR�AK5k�tZU�3"+&���u�� L�m��"���p�`����M�'|�ْ�+Ssx���[��u����U\.�z�����
���U��|m���PU��8gU�`��c�R�w�Z��� �l�g�`�bґ؍�y}H>�T�bVi����=�՝� Q� !]���?@T�>W�p�O�;�hzF/l�IAX�W�}r�n��%X&�o�M����\��,�HRB����=����[;�,��=�5
5t�N�ƍ�eU?f�XlxVHYEB    7744    1780�au�Lٷ�۟Q��na7���ζ���:���]��k�(}V�KN�R{�n��A��t�	�f�¬�t.I!�;i�
�m��Gɧu���A(1��𮇗1|��^��~m�|Ba4 �*�k�I�mE~��Uj,fD�wVK7�H5���(��PrE�|3�D�{���"#j��t?�N�� ��2ec�E7��t���yLY�l�c��gV0�5�,��
�Ij�b⏫ˎy⡄6�v��I-�Tgc��%�2���/�cU��|�u��Ҳ9�dH���~�3��R���:�p�M�N��:%�C�_	����$^����؊{>�x���4G�_J��ͼ�hANlq[!n\žP�fB�U�%���!�+�X!2�zO��ZF��&=ҖJ���]�iU����i�#���~�QM�;_^1��^������+�>��ac!�B2&�GG"��M��`~m�>\%� X^-h|P�E~�� �bIw%���+
z�:>N����"�ж��f�خ�֌.}��E+�߲V��P(�ps��3x�wPΏ�o"��?�%'�/ȥ[���AI=�25�W}h�K�T�W��톷�3�o�/�
�^u�.�6)��[@�_�R`ZW'LXf�uwv�aD��Bv��<�:���d`#⨜r�օb3�W�m_�wS��DaM�)Q�~<���;��@��xS%�lB���h^��*u� �v۬49_KP�ܸa�����!�������3�����c�����zu�=RV6P�&�:X�����H���y���.]��_@|�2y�CP�~b��Y�t�Z�7�U�Iev���b��ֽ�c^t���k]��.��i-<)e���s�A{�d1�0�L H�����J�J`lJyhp��T@��bJ6���zM�'�0�I'���n���I�^��D�ͮ��^LV@BQ���q͚����%U����9�P��rX�BS�c���I�<�7�����\�;�[�ۑ��j��8�vbȮy�|8�����>�hӊj��Aщ����9x�Di�Ի��T��c�ĭ%F�Ɓ��&!,gj��Zx�c��\L���sU�bސ,:5"�*�Ѳ{�Ğ[L�|��؞�en�;&�~�}��j���1������E.�w�w�US�����n�?�r�|�)ⶫm;�_�,[������<�
a�bѓR��՝K`�(^��ƓC��"N�FM�É����N�� ���k,��%��U�α�oib�ZNɏ[�@�A)��b�5�'֍��dzm�X� {5U�v��1͉3?��e#��U֜^����N�	=t���Q�ܿs�u����Nw�ڥ��b��cs�0����	8+�l��[����2	!�;L��V���]�ȿoi���n�Eǿ�H)��.��e`��7LS�k��X;p���L��
���4s�Y�'�,���-jI�oo�gB�i՟��2�y�y�x���Z��hJ�S=�o���ì^G�������K����*�L_'/T�ŚN���{mՓb����%��܆�+�qs(��5>�e`�HJ�,����Z������s�`U���*kD�1��U�r�쪘��o��%A��Hn�_B}�ч�<(6M+�����ngi8T�M�J�-1�׿�S�gdӳV�C;�tlEʇ���X�fƦ��Ir�E!O;ؙ<-��������h>�X�����5����Yg�J(WČ'D��(�tQ�8�������N*�`��7����%߿f�0�����ߌ����W��q�j�z��ˮ��*��>+��n�l5����#��?�p\3{=� ��~����^�ɒ+����xo�S��{;����ybs�2 �)��2 �O-��B5��@�Y���4����.Ÿ��\3������e�z(�)>��
�OP�ט��լ�҈h%$���AQRӯ)g��N�_k�~�q�[�v4��+�����/�еA�0 ��{A߾�O����sF�"���KX�������r�V1����~��2BO)�3��!K,��
���z�j0D��|4}/"�-��z&&y',���
\Ro.��1������_��.A��r�=�Q�ŵ��[ ��S& GL-3�)�hs4�?���{�*���;��y/�[�M��y���eW`�O�!�1vƬ�nA����i����RЫ������G���$��&��������cUKS�Gw��C��[W�t�՞���.�$�wkU��ോ�s3�m��-�!HE�ty�z�G�&��U�5Bz$�༹`����/� ث��L|mh #��-N��g5�HpLh���d�ґ�)���s�s��u	��F�Ή^%-��!`��>/�b��B˭�~A��*V��5�E��G4�I�����I9�WuRe�_�h��w������|Y|��ѣ^�h[ ��W�a9ũX�������q���M�A�w`��bA��c�B���j�Z�$�U��=�!��N�G���JTw0��B�k}�NהV7�gv棟�	j`�Σɻ����ޒV�ٖkԂ���W�y���d1�K�����kSep��+�3�������N;��26,���_ބ����%2:e���5��ޚ�o#u�j&?s-3N¸�X��f�0`���N�9���D����y��%EV�W�P	\�:W�9%2���64T���r&%2�F�C�ׅ���] I>'@��qW�s��zgh>;}�;�g+�sD��{�E3�ix1�8(�C/L\�����~"^����?��8��7Z��$��E�F^fV
��u冋eW��+�C��O�;�ڤЙ0��Œ�A��.|�+3i�l�$Y�?�S:2i�q�`rM4���Q����Q�vs��3���ymߊ�*La�c
�d+"�MmN��6b���)�a����X�H�p�t��EO�6��R�,�}&��\_o�!h���Y�͘����L����F�$�Cv���' �,r��,��v���?腧�	/Z0
I�I��%���BY߫�A�ѵ��-٫���#;���@ig� �t9��`+-[�Ubi��]�h���[��	�:�Sc�c�c�~�@5�p���O^t4���y��C�^�ϛ���?�;���\']�-���HP��^�� 5gƌ�B�o�ߞ��z���~c�Z/4o�zw"��>�s�()e���)p�e��#$���\ �a*�B-�����,��r5��@r"r��c����P�KJ�`�9������:������"����]�X
�jH?�;u�o���,��C]�N��[�)M�r=�$���j0�v\��#���E1�'5�X 'ה�|�S��ï�T��/������s��,�z���+���I]�%v(I@k�f��ݟ�z;w:&���Ւ�=��V�̫6�lro��D63�����L:����pM��E�:%�[V�
ο^�� {/^�6�]_?G�� 9�
f^�-i��� �[��R���9�36�b�ä�m\Oh*8�
�A�(k��v���� 1��\�h0d3@0K,��h�靈�8��U�V�vQ��<d�����<J/I�Ih7Կ�\D�,��y/
�x�<�苫���%��7'6����Ђ9����wK������ߤB?u�	Y���Q�|�aP�nJcv{��JQ/�K�zBc�FK���Z ���Tیg�3gGLy]+���_�(��ͤ�ƭ�m꼘�5���*ó���'�-1BF`E�&���x��g�]B�oJA�����\O+y�^�79A�$�u�m�6��{�٩�"Q����"���u*D2xM�9�ܷ9˜y,"�y:��B5�|��2����~� �l�����_py��Ӏx*H�%�/V{�e~d�䳹o*%"�`?٬xG�:��d�&[5` �F�2��(C�oKΥ��(o��-�Gً~�F���@Xؙ;/�P@;+�3��W m���G��+��	�"������?�&�%�[�h����z������H�E�k�R(S/a0]"�rpǧ7�e��9���DLqar%��vN|тaI�����|���,^�UY"����y|�k���J}0�-Y��!}���2ٗ+ڋ��?�Y�~x���])��X��b���=;��*��c�;��#	AU��P���䦎g	�ε�Ǌ��*�䘻v���
0!4�hU�6�#@A�mAf�i|5u��)%�,�e���b`��^���}�A'�ҳ+���̒,�K�EW�m�]醜I����3�,���Wl|��U�rl� �3���Ż�1/�dM�A�g�sy@V��K"7�_6�M@�p1�P�G�o,�}�sJ��O��Yӫmz%�j�:Eq�R&*�+w��J�;�(Z1���Wd~���K�ҨP �(H6 &y�1DI����37�rhCY�O���1�bZ���;x��v.�t�/Ѱ%�lAnĦ)�<f7�ņ;����q��
ζ�$ڿC?��4�t�u��g;�'KtJ)֩y���3Z���ղm��,Dz���CwZG�h3��<��2L�S�Y�p���x��6�/n�/�d��T$� S���3dE�Վ�U4r)�G]�rU�*a�@��c8�`��g�����Sh)���{��Okt�i+2?�ET�o�c>F̦�+�z�ܭ�JՒm����`[_�~��6�Y�w����5Iڇ�m�,�ڐH)2U���K�Q� Ylrŭ�]����D8��h/���� ��kپ?Nt=����
�̪��:H`�>�x������L�.C��W}��k� s-������L	��6���^��[g���p���Ͷ|���7DHÒX�f�~;�DESR�iγ������
��u�_I�˛6�g�ؽ�� �@�P��f��*�<9V�V��K>��1F����
͈�L�#`��&�TJ�	���y� �95��sx��S0y���=d�}݂�&�9]J��%��yM����N�y}JN1)&���:^N��=�� ����Q��k ��4�ڮ0�D
⼉�U]"a%V�	��Yy~�i�ew������W��>���̊:"����]�.�ZLj�D0��������o��:�[�yĪ��Ԟ��k�u�u�d}����#F�, � 5�4)�D
")��i�������z�W�j��S-��K|�o���M����e삪j�Nሞ�N(bN�S4m����)g=B	gjd���jus�S�*��a[������y(�z���x5��$l������?���g�u(*Fyſ����ReE����=a�i�@� �ud/��k�"+�X|��&A��C����)�A��,W6'��eNW���o � �������$Z�R��iB�B� �ӺEEY���j`��QHp��F��36�njY�w%��Xdyu�I�o���8�HΜ�2��gK���Z�2�0����$e���; �[#�@Y�~��~\��+�h�vQg�	�\8Ě�B��O=�xp�� �c�k�Q׊�؎A?q�WڪDT`G��{�\#���z�Ѭ��5���oAt-��1����N:NL1��\k��9��=D�����5�^��T���5���`�#��zc��|	������������l�n̵�i��T ����΃ƠZm�e���*?��1I��-�c�&�����(���.�%��=Zm�$������'�{"A�4V��L4�9���	��=������^s�Q��m�����)Es:�����E�oFt�L�چ��6fv�K7�#�:���1�Ş�0к���m⟧��EVe��c�:��T\��,���j�DB��$`0�$�ܯq�
���Zo�go*��w��@l��q�rѹ/H$���t��m����$@����eD��Ƽ�s�|�pj�-��u���B�+��\F�6ۤF�P�MZX�1�_�e[�h�H�TB܉