XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������Y���Z]q�X~�����n���\W	R�@$��7���ֺ ��_���ZA&xH?%Y�r�&"@d#�%���U!�������_,B(�U6��4�޿�f�OY+���왠�^"*�,(�>`° �2�?��-n�*���sh<HGQ��N��F�n�t�׎2ƚ��.-��}2�f���̡տ=�fN�m��i�����JSt*:���0Omz�be���e괧�D&~y��α�봐]u�݇g ��G���A���n�XԳ��A���зc�Ȩi�c���w3�wuj>`_&�"�hU�eY����\K.�^���;~���yq|�g�� �Ne9�VVaU��ӛ{s��Dfp/�X�9���Y��C����/���Ft� ��x��zB�_�{�ۥ-�W��Co8�[kH�(u���M�����Ē�v"<P8���bf��\�8�^p��F�jЏ��x�
|���prJs��>������J������&�>�8�Kg�' ',Ty�ұ�7��� R_
�C^��Y���#�����	R�!;�h�Ϡ�c�F�/N>נ 
>|�����#����Vx�%�o�?`#n���:-@��{�B&Ʌ����õi[��~;h��1"2[ɪ�k1��n�j+}����U!����ao�F�4
�C�7V筏F���6�8wѻB�G ¯���>�
�r	�N�M˚AJQ��9��s|�1����ňmW��_����XlxVHYEB    c763    26003��������.�.���~d�J.	ZY��ބ�mӣ�Z���9f�S��n�������'�>X��R���A)кS���OG�]ԋ���"Ý��w�+��o�(`t�7݅�W����X�N	$Z�Zux�x�.��CY���=�m�2:-�$��R&��˴�wxu�$�>V/�R��چ��^a�@L�F�B���P��]�/�˖@g��q'd�]JT�GM!Ws�,O1�	J��sFV1�^��"%�eݖ��:)uWu�m�J=��g�.9��DJ�r��%i�hm�v��v�B��:�\4�lb���
�����0w��)6*ć�FЪoO6��a�O�@"�M�vR+��9��qrv3)�ģ�l�k�t��(8�2�� .a�-`�jbe�-pr�V�5��%J}`w��	£�F=ɀ��Mp-��t9�L���}�W�!G��3.UD�z��>��_ּ� �[���9I�'&�G�[N+����Es����3Z���T�>�!|�4(�?2�Ń��������Ò����C�b��}�4����KػT�o�4����ȷ��ݕ��S��Z��a�0ִR��:"N ��zNߺe<��/��r}2���,�z�6�9�m6�=���h�|c�M;��n�30�`?��R4��6o4��F�R,�D�w[%��|���uл"L�N����2��T�� ����� ��#V�;͑v�떨q���BI/y��xh��"�E�#-r��L�`HV�E�<Fq���ӌ�v�!���</*����<��Q.��\/�n#ߚ�@ZU�m4qDʄ�Az��4�n�:,��9��R*8�7i)��=B��E����0=�r�����za]����g�����	��"����b:��.�	�s��"Nv����v�C��ew�ʁ�7璉��v~�ϤO���?��w�A���mWˎ���/$�aߒ; c!>�&����
��K�1,Rk���y�9(��`���������hCC�hTmHs�+a]�DCԪh��k��ɞ@]f~�b����}��`a�z�噾0�@Wöd� ����e/�J��*���n����(�x�HJީ�_�����E�ݦdB�:���/
�X�0X,��^��i��|@ �Y�,�pzV���eX�pm�D	���l؟PV�O�@�ŗ�<
�&||�Cd'^�J�E���jp�C�M��O�^�'�xL�ش��== �{�d����Fl#*�;�E�k���l����[�È8d���K�JZ䗳�t�$s��x0�Z�o��w)n(	�'Gg�M���C���z��
�~�|4���bw�	p�mp�)����/�"�%�y��JzЬ��QM|��T�쀝�%=yK�5g��Rrz�I��"�UMOO�bD��|��h&��lP���k�&��S/qVQq����vc��ɜ#/��z>�װhz��?5p.��X�fA��~"_3�N`�De�̢��$��Rp�zl�V����	�����&��+\TYW{�Q�.���/NH ��Kj�ҋ=<�Ѿ��&5�L����2�=��t48/�L�^F��n���R��y��}���'0��ņ!^RF^uq�զ�H�8�R���O܎�:��U��R�RB�kfoi�'��
V�Ⱥ��5�l�KY�0h���h�<@*�ե��]�@T4&�8p��G9��Vb3V���H �������۫�<�*ٔ�G8�=����Z܅<%=�a�9��x�׉O�̀��X`�X�>��������~�31=~�G!�y��f�����z�m_�!�q��x+q��(ir���u��P4DḰ���!Eu'V��kY�Ҡ� \��C�\��&t�����I�)Jfx'�����Z�S���o񎄢x	�狓��?�z<;e����;_z�/gp���#{h�7��f���(Нu�4G_c�It]���있Vڬ��.^��N�t�wn7駥?�J\�|u�g"6AY���Pخ����Lr�db�@�?8�a@�P�@�n_U��M�Kd� �DE3�S�ky��6t�D}7�>���U;�v��������������ld���%���Dt��8�[<C�G������%�p�䡋A�u�g�\�a����r�q#��|9i��Fs��a�ة�	��P��몣�	jڳzA�b:G�KK���
�&����F'��W�>�wef[4"�(W�̷��{�����(r����[��ͪV����I�xl�//V$�`�nq<�H6�@�;s�v�bd�M�:7�2�:C�P?�C�3��t���$]=V���Zt��4abh+�=�w���F�I�F�f����;UTC��j�q$�
�'�f��k[.e�K!�#~���.�,VMԚBl�yx>\�����|��D�����X�7�re\
B|���'��'���J* 6m�h�?%!��(I�e����|��;/ S���m!���ä�۸������?�K\�Mso�fU�༿�f��[Þ���4�!JU9�8�gpH�^u��>�b춯���IO�[�J�FF�?Y�n��R���*#6h��|Z��ǵ�J��O����āw`8����XٜY(����)���ڲ��c�����=l�V��t�Ŝpf�VmŖ�")��RF#�O��,d@h\�4�0�u%�!��̎\ ��I�u���F-N!^Kc9��d���1�\�|���P�4Z`iF���J���V����(%AU�D($�c�o��B:>H8��e�<�a 0�o�Lq��W�wސe�9�����>ua����d(��l�C�̊c^�A,�zҷ��E���H=/ &`�v��z���$-Y��:c8W�P�r���t�1ì�f�\w+��-A7�[WO��\��J�N��B�#�4û.h���p�����W!�Cy�*
�=����FY����>�u�s��FW���.b�
4i�4�2�A�~� '���Zy�B��;t^��IKX,٪\�4�2��*.���Wb�Xi���>��T��륡�O8"��Z3F�6��T��o���Sj܄�ɑ�A��U8D��}Zu 򦏫p0�L#��m+��
A��m�m9�?�ɝ�t�!�5K0�^X�V�\��� W
��:^�����%ʡ!U	��ݦ�is?������݋��C2��p���/���~N���j
�t�+	��*9���xG�O!`j��'u!��|	,p��G��^��_�o��1�x,����ASf�6������ �b[��ɰ�a2F�_��>�#��C����)x:]f�1&Գg�:�k������R�ҋIq�*N���u,Pq��Q[a�(�d.X��|c����^13b򢝯���/@�28���B�,��fpN/u�{�a�5�"�5�}�@����"K��N�4��:�3�|�֎�	�m{zY�P(���G�H��>M��z�����E�a�Z�
<�*��kp�����*]��c�kuf���9S[�X�m���аS���I7����=��T���N�C{YJ��y���ᗽ���t=��H��;�P}�Ge�����["�JI<�AU`x�1$ܕP�^�f���f�]<������3�̝�+�������!ׂ}�������v��v�q⡞�/Lr_�m�t�4���?����R5�ޗ&/ҏ�������ۉ�Vf*�'��aP�uZ�U<�������ՔWoT�^iC�?fb�|�^��z=�	�rc[���+��"�IMV�c��8g����-bC\o����{�-� &�:`N'|ϲ�I'P��U�+��u�=�0�=~b�ҝ�ҧ�X�7�#�,��2�9!??�H�.���Q5��2�uLwG8�nY{�:��9���a���jJi�0L����!�0y����	F�'��l���)�`���bi���\Ѻq�td���W�c�]p�︗�hh�ː�J���٥�w����D'�.`Q��~�ᒸ��p�T�3x�k~�"��PF��@Ks�����41�ݢ�C"@���&m�r���T>I:%wtєx8�/���ISu�צ�Aĵ锌�8$������|�9����dǺh��ٹ�5���s�5[�F&'Y�E�w�"�\�������4�����Q�)Y-�,�dn�䅩�D'�[��˷]��l饰E��/����C�җ'�������?�Y��[�3Tk�*neV<
����V�ӑ�f�Uܩ{��N�8�:��\�vʀ-B�<V?�W%����ы�Z��H����?���DDTJhÂ\8�� &o��x�i�vLw��6���x�HM���!���~��� �+l�9�
?��9���o��tp3uf9���D�gm_?Y��8��6R��>px*j�;k|W�/��Z�q%2B�r�)�(ۈ<�e?z��	��J�{Ũ�2�{�P|~`G��7z�;���T�VqT:�Y,�����N3~�����
-R�!,{�ϸ������!^����Aގ����T�"�gk^��s��O��߀�E%>�bŎ0Ep^�vw������s�$�&�]����ww��+��9����*M�ʖ��hhP.�̦����I3zm6�U�#���!����U^ż�+X��;��1����{�m��RJ��rAo�zoR�a�N;'�}�z�v(4O�>�������ٿ����y�uۭ;���b�1�S<E�`��e�P�\�ձ���jf��<������^�5k�H��yZk��!�Y:���B�n�綜+
=��^�,Z�m�Ȓ1=�e��8�hu��o��۽^Ş�y0PS}}J���q9�ʧ/0�ʝ�I��	�x*p�V�
�24$�a��-BS���C>rz$I�p�̼C		������e۰(Sy�n��FfYD�_��&��tC��&�qf%O��|��)���*�M���2R�J�1/&��!X�hgTy`<i�-x��R�w���L��9���h �P}1?<6U��Y2��J�f��⏻a�(RX�g���O�t�&�̵W�����]n�giou��t@}�NZ�!�C�2#�?��x�����Z�bFQZ�ꟸ��)�3g���d��$C��p.��޼��<yq�er�aQՔI���;���4���@�'���	�-0�����9@ly9�	Q>}pEv�O&bF��j�D(���کA���q;b�rw��)�!��c"p�?&���A�]T-���l��HI�lD;�<\��!�	t��Q
���!y9�6�і%�)�ާl�2���<��9��n�ؑ���/S����I�ô��	�Ö�]Y���,)$���������N��/A�츕L+�0㯻�n�� �^��H��U@�֌�J�-�FY�R~���G���*�f��;΄��\�F��)��a�� ��1�[�ձ�{%\d$]8��Q�ݨ	�nl�xK�z6Z�-0�����	o���xz��d]����3U_{0���9����{�q�AY�2�^xP�@�gSoߎ�9ڈ����9�i��zrR� ���f��zA�yO%����1�ݮ3�w��]о�o�Z��!>b��G~�_~CT����,��D@�� s�r�[Z]��g 0$Bb�yǖ�8-���a��W�"�
����|j��p�L<�[j��Կ����kX��3C��n������tR��-s���Ԯ��a2��Ԍ>k'�t{���^���t�cg��/���6ahp��ZZ�i�P-�V��I��%�s���I��w�vMϝ(2��x|�%�a�z_i����{�D�5B9�kgM�P%Z�@��#��s�mi�S;bjŖv���$ �$Ԝȵ��Nɋ�A�P}���d�v��&����|,���C�S]s	��ӡe�����c
{ǈa(Xl��,�_����G�ե�C��դ�\��Ӷ�Ng+��B+���s���2Q4�BG��/��x�j�[Z���ݹҫc��l�Lm+qYg�������+��hf�4��=�UŜ�4v;$~;G�-��ҫh���<r����'J}4��2Lo��M���l��U���+Y��v4�ٻ�a���[4hh�z�w�F0��c�g�Z��uƽ��D�-9v(�e��4���3��wPY�C��v*,�Ss:��f��:N`��dM�(�
"NX"��r�X���u��>4bs���f$�E�e- #S��}%_�n�C��ol�2��ĕ[a��n�l�w�nQ��%�LO&�#J�	�u^����i��X�qz�S\�k��FA�`m����u����X#c |)?Bd������-�O`��k�py�W�a���~��ΎA��/�['�e뮠�Y�:��rec�:���Oٌ���R�B5�_l����'�d"ܐ;���r����x(uN@��S�e�*]>� �������~y���WSE�l3�%�vY+���ն��Lh�m�ܡ�	��gIFup,��>$����v�suc�9��=昸�L�����D�U7����!R��醣��_�;J��J��{��a1�ߙ� ������(�uL�����4^V@�|�Q)��GQ@c7�5�Ap�~,���	hh��{~��^��*3��ݻ���l�)t��*��
�p�H�����dqe;Hq���)�Y����؈���r�fj��xլ�*r���ʹ�i2���!������}�Ed�{��-|�\9PT��}1qG�~4H�e{���,[Qb}�{���3���/�ՈUÏKXs�jⲼ���4�ΈVQ��>�t%�q�G|҈n��gx���`:�^@H0e���*�\[ Mo� Q'�dR}?v,�m�6Av��\�oD&ۦ�+B�9���U*�@Y'�<Fu0��0U[���mk�t|�%12��<�I.u\��2�U`^�3Nj�TX�/�ѽJ��=�9�PU�c)E���ϴ�g{l����Գ�y�$�	9󜘃r�2��kAz�s�Q�Q#��t�$��"�o��m� T��s�T��Z"���O�o�E��4-���4�._���t�4���2���b�Ŧa�u�W��������Z4�^�w!l�#螋C���ģ��sX/�E�L3�'	�ގ�Щ�h��oU��`�br��k"�i�74H�,�i�V�o#GU��/��2������>^�览��_N��δ��b�jh��S�i�U��o�#R��+���!��h^9�D�T��8��N��/�th]m��M��L�o:�G4�n�)����vLH@���Ӄ%�x��O�/�[��Z:��<`���=\�<긵��J���u1��Z�����}�kU,X��=]���1#�V�(��;q�'Y��B��=K��d,��l�xM|q�U��4��Njہɖ��W��r֧+�L���S��Y��}�@i�A�j�(=�����6�����z[��?ZD�[�`f�I\ 5's�s���?������#�Vՠ�C�~y�`mci¶���KO�0Ƈ.�_��\�����ٞ�~{[��&��1��^��@І�	�Hc]^8%������7C�'�39�&��������'�z-:\�y���ם�Q��m�T�j%4LΜʭ3M9��k�W���[�@~Ȑ�&>�R������GYH����w[ޜ]h��`�}�/0"����	��ں�{�6aГ���}��%�9��N�R*#_t�9�D:K���l�ϋyW�y^U��"�k���W
�����"�li8C���wB��'�/�6���ݭ�х�5c����Y�tB=da�D�E�$I��J�˪j���t�;u�����xbR\��/��JB�+*�͙?����]ȎZg�TR��P06����*)��p��|$lQ�LB�mк	f���B������%�r����s!����h�"t�xT�u;�ػK.薶Ofl�6��aⓋ'�۾y�q�����I�������u�܂�3��9��D(�HQ�	�����g ,)(��p����D��m+8^%�BO��G�	ކ:���	�܎�I	����HUC���zF��H�To��D�jΖ�@�[܅���Y�j~*�7����b�$'�1ŹI:���cl����[��2�$�?��!�����U�E��j���2�f��i��(�l�����I�n�7Ocs�|t��=��/@�jڌ������[+�#���[�`���m�a^���=�J�3mO߼��<�#l���)(�|!�j��g4���Hi�pQ��3*Un�rv�yj��ӌ�>3<�Ω�y6�?Mek�:��� i00�]�Ռ|ɘZ{�+��[�wV�l�$
�B���&,h�70de��ʙ
�
z�d���&��jR8uN6�)¤3���S���q?)�	�>�0���I��@'L��E$H8� �ړ	��$G�t/9�W�0�Z���7�@���{�g���X��l�����3�WG�h5���d�t�����O*<��\�2q�t�"%��O�x��v͜�	���HO���@��׵��#��}K>���b�w��EϢ����rNVn�ݘ_�l��˾��2��t�Y�weӭR�q[�L��,�� ��07��}SXC=ԋ��ҵ0�4��ˣ�X��?m��G�F�/u����š�yo��ĕ<�u4�N}��̙��Oso��"$j�L�2� �'sүk�߅���ϞP&U��MG}I�g��g�,#:�B�>��y�|�:�(e��P�xc���� {����I��]X��α��(��
����\���&b��1V�E�`�A��ǣl���F���g��r�����Fµ���̙�赢�k�]߭\�âz&|�~�<=�إ�U��= ���������7d��w'��F8�K����P�0o(W������R����ɗp���+���eg��c� �l{q�e���x�(}E�v�_�j�RT�+���d`	�~i�=�'��'�3)�8��`�HD��Gi����&�U���l��;����E['K.N��w ���H���O��	BA H�u�5���_�ɼ!˘oBӫ��A���c�Ƚ���.�P�㋑bC���1_��F��a�FҎU��_u�Q�v9�G��;���`~��� ��l����Q�H�w��_ݨ��k�N`�ң�kXw��~�Δm3�ҭl0��LA�F��a"��g���t� M~�"�$�5�T���1�cƼ��B��D�j��LŶ!娣�XU�h��(��nN��~�����W�����x�3���e%m�
֮����p���
��/��H����*���� <w�
��ډ�y
��I[s )��G��E�d	 剦r���yKj2���H5����N��`(E�'M�G,2��LקV�GNO.��E�p��@��a]a{�_2��3��}�+=�,kP�vXD�=�R&���w�ue����)�Sb�f)��������|�m9@cXޡ���?Ӵ\"oQ�� a��N�^�
(B�y�bͲ�2�z�U��2�/�[��EEbGV�B�o�|z}�
�0n]�ٸC�I���'�s7<0�>�Y�9m\Q=N�Њx0\���mo&
1PMo_Ƅ�O}u�������uт��