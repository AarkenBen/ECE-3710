XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��Ͻ^���̣��_Q��I������=��Mg�*�$6�;�B0娅��d�O�-�5#�hZ�5��t��%5^����
+��r���������z�e���$g�֭���rp��q�5C���Q6z�k�O�Wϔ�C�	�Y^����Ba��I~&�y�����>�ʶk�`%F_�MGӫV�M�r��>=(0s�����Jo�2�o�(��9lP?_`�&}؆�iK�o�ԇT}ˀ���c�U�'I�̤�N���=q� 
lQ-�}.�e��=�����"�Z�wBϊ���C	Yqe(���v��}<�[�ݠ}?�n�jblJ�5���P��<i�N�u��P9F���TJ�id�W32!v? �|�(z�����`�?�j�K�Θr�دW���(8Cjکg1�jĘ�Q�����u�@�^���RBw�?��6��v"p���V!l��/�r�UIv>��m��;��ŭn���nl(��>}�7W�x���ŉbZ��/k�$���#�u�|��Y.4�49�e�[h��$��Beb%��mL9�$hr��:1��"�������]�*1���/^�YX�k3�������L�y��3��=�66�(`�I6*/�~$�+�	W'*R~���C�T���߆����_`o ��o%��.�8�8�����Zl�=(+�$���VU4�v��!3#B�X��3�:�D/.5��h�y@�F�z5�(�&C2����:f��li��Z^�hQ{�*��XlxVHYEB    aa52    13d0M��&e�;�7~����>Cb��1@Z@�Co���������f��b���i���)�0V63puU��6��S� ��=l)CĽ�t����������NQy�ɢ��e2�g2e�ʚ�|�8���0�"<_d6����k_����7]:�o׺���߫��V}~ʗ�B�]+��?1�7�����KU���u��g�!�6���dHl
��B��H���%�>� �� ZF�L��VN��Ɏ��]�
�\ӈ^�Vg��'����v�����C-��)���'�#�dAN��]Oځ�/6	h���A��N�`�c� ~�w�qJ ����|�-���z�g�>7�36��!�ɍ��|P�]#�E�Y�D$��`��"�-�/�	�Z~Q��Z9��ee!=��\y�]�E�7 ��޻7������M\�H�����{F�!��|*~�&ag'��ь=��+|`y�/пQ��PѸGQ��|���3�`���eYA9����v%kv�p3k�ycے�Wt�e�mg�$��N��� I��Ӏ,�.F)ۯ��e�΢��C������tkP�}���/�)�n����y8�]�,�͢��uK|)��u�J�QT����܌�VY%� �f1�+[��Q�ӡ2S�P�@޸D���GXgL� ��ʑ��*��,|���u�8��ێb�a��z�?) [����.ߝuڎ
G�
F�W)���⣻��k^��$a�p(�X2K)Ќ2a,'X��?�)BH���h"�z�-�0�W+MA0�3�����[Ǔ:��T�^-Wt�{� `�W��3�Lq�f�eUbkg����N��\:���C�-�Rw���2��H���n:m��	�����;��k�j�������Є�<5sk�A`潨�KB������ʍm�  1����a��PAM�;����0� ��B�Ý�P�!���f_[LWt��H���'�Uf�������;�P��{�a	9����+��??C��GO����b�ta�f&n�2�E4
���Fa�A~�v�F¿/Km�,����0x�f ��AE{#Z�}�Zxƻ���\!	���R���t-kDSs���D�+�	0tOf�n@�sP���VI�'�	c�&ӎ��_%@ OGô��_}ӵ��?�dA�_��/����-Ƃ`�<�Ӹ[��dԫ���h;���p��+Ww�e�C`�0��C��/oa��V���%�rE��I����1�
�`29�$޶s����m���<̒����f舉��� Q���8���GύWI�(����X��2xO�h���A�nh7��9�y�E��&�Ǯ�hT��q�]��p��y�{��LAz����Ź.�'WO��������^�s���a�=�}5�[��A�4h��KmE~d�
M�'>���2i�2�n��n��l�	�ڽKC����}�k�7&5j�X�D���4rƐQ��+5�����i�@*x�'9	_.M�M�e��D�� �v'�MxH�]�xX �T��E,���>S0�o���qi�iʅHU�S\&���[�HQ�����i�ɮzŠ�֎�f��^�U�ma�s�wS&���4�燣������z�+�m^|O� 2�߸�[Xǘ���~3�c�1$�@s,�ӊq+_��<1p�[�����,�g�� ����e{V��9�̲b�( 2�TA�*֩�4\ӟ툲��.&2Йr��6O���7��Q́/�:��>�������#~H;�)�|ֆ�ѫ�zԿ�M�В5���s&ūo:=�<ۢ���u2��Ý�m}���!��!�G�'�jviox���k����t���p�����q�k��F��ik�|�[Q�q�@H��L)@���a����e�.�Y[�X���Q���u�j���C�E�ŽU�X������&A��FaU�o^n����ș�)P��|�c�	G�nAH�����D`s�tV�Y��T'���B�X��sn��̡����Ǆ�a�rʅjd�c(����vH�B×�9LI�kx��dW�~e�������%�`0ȍG���P�������J���)�;��#�/�V�K�-DF<%w�>����t�W�[i9��vss�&E0{�� c���&���x����Y�������pZ�_�������o̪�r �H�+Z-1
��� ��b��c�j����pLʁ�#��Ԏ�U;k	�E̿��B����e� ��Gƀ� �$�SJAI�A�
���9#�"nd�Re�<�̫�Ԯh���@�P!�Π+�BW,�� �=�Q�+~�nM�%�i�4��-�|"�vטz�<�rf"H��+c�^v0ʽ�0d�]�����<�^����Np 0q����T������5]pƄiu!<+���<����h�^���I�i#�N�q��]>�EܸH˧`���~�!DU�����_P��g�?�m�&�✵ϔ[[e��;�o��EMr&a�;��؏�P܆s-ݩ�������u�y_�DE�<ޖ,i�:k�z��Um	�{��F�����҇Vr6<&%3������؀@[E����G�y�i#�����b�d��WCdU:n�N%;y4r�W]�}E�[.)&^����;v�n��Y�IbtzT��3+�� ��_�7��%���m��te/��C��:N��"A�/q������ȃ�KO,�*��(_��',-9�ӂi�w���.U����f�H��"/�1(��| ��ҵEn�|�ОѨ6%NK���jx��ŋ.�e��\k(-E�z����aс��X�v�n�*DH� �I�zN\�:N~E�}*�KX�Z0�@�Îo�#ߑt�{��?�IK�fV�o$إ�4 ��=�;9]�A��R>*���?4�z��3	�?F�N��;+��e�>�Ǎ�� QR�Iƒ�s�DO����d\�N�Zn"@H�;�틎��{�R�Oږ�"��a������Q���Y`Q�R
���1�sZ����3G�y�\� (9>?v���>.�,9�|��7Q��5�ð�ezK(�1@L� ���d��s4�_&�)N\Vf���7����  �B(����W���ueVt.Չ �_ߜ���p>��Z�}E��	&p.ե��y���=���:�g"E����E�^�f�*@�0����uZ�� �%{A�W���J���ֳ�ՂW��*"�3B!��=�
�CS��5>gg�L�x����-魈��ȖvDmB�w�������GF)���W:�gR�q�3!R���<̳�C�v���zS��w�;�6�=�.R�^0c��[���M�n��KT����<�R��	�I�]��Y*����i�Rq�����\7�4�>'�c ��K�wП�q��8vK�04(�q�,XGp����PD{����¸��[8������NŻb��h��	̊z�f�/U�q�P�t�޾9�`�Q�f����z�b��_ p�wv:�F��W����o]|��ʕL�1+�{����?I��i��4�F���7_Db!5��P����T��P�I�n:��ûN���A�:�ksS�фl;�Sc�-���v-�x�y>��$k�ȡJ)�y8���0Z�u5�Ц����k���*Э�����w���m�h$�	�q�����_h����?�Ȭdj����up�^/U@������ǘ��fpФ8ͱP���]߲����J� ��;�H�Rd*"������T��Z*������x8
��	�d��$�����DHZR�s�5��ﮟq+�JG�NW�@�
+%Y{����K�O�A{���x������wu��;Z����[�n&>����?^�̙�|��鉾%����-�J�7�*_�cW�e6=��X@��\�4��"=<󠫑H��YmP�ʘ�7�������UN�����N�nl-�~�/?���w��)
���я�f�g��`R��@�aIG}���/=5Zu
��M�+;J*FG���f9��S�1{���Ʒ��.�H��发��!����A�@S�?E�t�=�3d�T�$r<eˡ=��^ ����L��^P9�WpD|� @餕�'�׸�K#��/?���H��<L��!E��_%�n��kn4�4	��0�Lp�wU�zzeZ����G2��3�*̝�䂿^-�7zx`C)��U8�N�a)�:&�b��cy��_[���x�^	���>fn��+Ir�^c��0P�+�[�	%�/Q�q�-'/ƭI��C{�:�f>oG�=��QI8OS��sR2��b�.Ґ������N5���PGLh����3��@0�2ä��xL��5S��ƖN�VN1{~�ٽ%��ʽ����Cd��]n�E�v�{��D�?�P����%�>+�Z��Ϡ.敷@E�8w ����vHm��޲��XBU�,���>!N�r���V����D��V����T5���<q��Z<���E�>�b����C�������љ�{T��]�ګ�+EӋ�[�>\Gz|ӱYp_I_G�LN'�h 9_�(M�q���H�4�A�����O��k>H�_�l��Y��Z8lNWA������H�ʦP�A O��
!����[���[c��V�ҤV�3��N��7��Vh�T�E�m&v|x���p%9�0&�F�9�Ҝq�t��%�t�X���0�g~����p�Iu?s�ؠ_�@���ᵣ�s_���S��{G�f�� ��Z��r�w�2�����
SNǩ<�I�=U�9�_�ԷG[�S��.��w����VVs��[��7�
�w��Y�U��v�p6����X��U��]�K�б���������m�B*�
m;'L�]�٠����ʤ�^��\�{�u%�-������6A[��n<��s��_<�M�&�в��T�^i�I;��B"�Prh������t���W�G�4���\�NV� �@G���)9��8�D4X��Nx۴���!����8'����U�����@�?gX�V�m��6�a�����Oz�ˈ��J�