XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��=�)'bn4�Ǘѭ�j?;s�8�#�A�i��wy�/�7$x�����7<���bs����?3���� ��P���&���k�����e� �b���0�I��{H�ݤ��o�=�ش�}��0tع���|�Qb�1��l�¦�s��Wƾ!ŷ$��L��z���U���*�_�}%�U�=V��v�ZNq_�93�ަ�xq��W�(|�I������Y��`g���ܑ0y#��%j5�q�~4z��D+Py���f���rpS���P\��׃�L�֝Tˉ/�9 ͶS�n��YF{^nr�}���RJ�"j�\��̈́�}a�h=*�߽���2x_͹�6g�?��� ͙�o�w�4����)a��E�jVWҢ�/��YH.w�O��4��zI�P���ݺ�B�2wJ��R����G��$�'��i(_6�7_=�v��w��	���L]�5�˞T/���!A���lV��D^�ή�T�˱c�ao�u0+Ќ�J�j\�f��v�y��=����.�+��1���}g���Z�+���oԂiȍ�j�K~��l��f�:DI�������c�W�o���X�+���3yQ���S��sU�����<�����d[�h�,Y��	��H��N�HGT.&`�|��)�,����2�`��7���Q��o����IB'O�-|��+��(�mO܄��7q��b9<���`=�p������ڰ������Qh��3����U�s
��+x�Y���u�ga��+XlxVHYEB    fa00    1790n�P��;� �QJ]}��[i�m*-�}�?
���5I��Z�D�N��v�\$������@���F���db)h���.ď�y�N?\5A��zw�;3'l�}(��ƅ�P��際�JQA�ow&��Y�����^"��l��Y���i�Jd�Ր�FH��4��F���/p���$�oA��F���W�#�%�V׹w�I�uO'��U��1_�)���R�&�?�Hk�����a��!�G�`���iʊC�|M(����>�w_�C:K��dp&�ή,�նog%�Q������ƿ����-W�+ai{E��v%����,�hJ��BL�
��=�H����H���0�\��^L��Sr���hBUn{��ZW�Ъm8�i�:������)�-�������L?[ꏠj�F�L�^)�[�%�9oU���N�d���6���U���!�,A�����p�w������'����	����}�?	 �?�0���m������'�Y��T�\�k"�o$\��۠a����5�'���=����`�ו����ޡeظ'd'���q��E�(N�/U'��p� �khB�%LKx֝���'�����A�'���DJ##D��j�'��|�ہ�\��r=Hc�����M����A�S,��;���;�����AM�R`�-���4�j�u3��l[�?��kr���D�ɓq)�˓߅��F��X�x�S0����H�ԑ��)�u��p�S}(�_��&CRE~i+&M@�q��>�z6�(�M۷A�-G�'< �Ԯ�
����h�v���+�س�|�4)��N(���RvnC��Qf��dĨ��NP�*��d
��{L���sQ��"��`(O�A��j\Dx�t�婛{�Lu|�JݻW�q���%׋'�ޱN�Y� b;�7��3h4���gW(5�w�!��;�(o6cN)����љR�X�|D@����}l-�"�E�b���|a�Lz�A�Ҁ�	�Ls�
�C [�)��i��T���[��:͂��ID��U6:��ӵSJPwX�{�#�}����CL��V��Qt�;�d�N:<�E#�ј+���	�C�MF�h��U���`�0B�q5����u�<A��ol��;�f��{�8�g_]�wv#��t������R�\+��_^�D���8'7����8�y�k�]<Z�7���>�s^Iγ��0�p��G��_ltu��3r�y7�R��kt���ZgS�*�j�SA6��@|���L"�È<'S�Ż�͒8�a�X�ߛ|r��w�`Z���Һ��>�;X�ئ�x�km�,�?���#W�[���M��� a��1�  [����Y��N5k�i1�5��7�z,��狈A$��zI��7�>-m�yB�gR%������[� �<���&fq�(�֎[;�u��rk-�#l}�M���K����S������|�|��Q��m��ь~�D��?�ۏR�k��&��ZK��P�]@=[�����"�S(�po�6'��|y�6+-{3�JR����^���&�*X�^v���s�6<�Ó�~�v�}���л���eT`�%Z^��g�Ԗ�+�M�u�^Z/��(:!,���g5F*1���,�L3���K��s'�1r�}YKx) �j�;z���1T�i�3(\|ִW����kӵ������@�:�rT�$_�`Ƚ�	��|��g_��K�1\��_��y�w�=���Z��j��fA�"�M�ۥi��
���pWUo}�x$xg%ԃJ��^�����mƦB؎��l�n]5��Q����x�������6s����еyӹ(4%<��t�/U���)��q]��+�ǔ{��fVOy}s��'/H��>�t���a�\�~oW�7G,$b�W	��*�hc�^۰	���}�yڠ�4ߙUr�A��Ro����I����~[9!�	Rqpb5)���ZxJ!��R������\U���_�1p�Ґ��P��B�nK�D���X��pr�Ke��=����5$C�b�n��r��?@#���/}�R+�kΎȲk��Q�x�ӷ�x&����!�Ţ�O�����S�j��	�n����w�����971͎M��C���� �� 2o��?,���MA�=�{,�OZ��I�:�7ظ���#�a�J�b�I��M���pK�	�y;ob�?�DQ�����G��5�j�ʫ �"AN�QxB�����c�w��h���K,��N��㍬�jڡtul������\9k�&7ݟK-�(hD��=�N��!Pp�A{k��y#F�)J%�F��Vi�=�qU̯���F/I�Z}����w���������xճQ���C~\*�"��1�wN������7�OD�߯�{���س�p�s(���K�~��4aj� `a����L��-���!O%�.~;��XMA`����i��}1�ȱ��:8��Ŵ��x<���&���w���?���o�5�/?��i�o���%��'�،;wA��oĠ��N�ۏ���=�Ǯ����⁙�ie�l�L~].X� �r���� �Dy}v:V������iU�R�.]ʰJo�����[@ܴ g3��D�ז��+FuO�S�PDY�Add�=��c��?xK���;��73��_ٱە�!\�xsM�����^P�Z��ԙ�/���߆�De����!�Ҧ�G=�4���1Ct�ng͠W[�ʎ�]���Y ����U�
Yn�O�n7[���F�	\��_.���s���/�3Q������'��%sP��Ԗ<�kDv_��g[��a�����r$H�.�Ñ
3��plwl�)�ѰC�3F�L���m[����tqFT�Ӈ/KV��W��������7@�l����bvT�xjP)z�����:��B�\��U�q�{A��7�V]�7�,�X�۹���_��Ju���9��y�mͳA�d,�< 8U��-�뮝�S��@�Yx=���˯���j�}��.��N�ko��|9��,]�N�id���(2����������,/�� �}:�f�ӧ0��Q�^����:v�B1�s��`� (x˽��
;-�x�?�quU�����+�<����4������Q�lp<VpFȋ�j�'�=�4X;�7�dƦ�� �wJT%�T��������� k��C��%���ց���#%u�`�wьh�Fn�>���[��~��sǾ�ː�Y����Ʒ�#��5��
�M�� wF�U�F׬�c溉�0L����w�	=k��}�le��JD����"��%�կ����ǚ��>ƀΫ�B	�Fg���ela�?��.������� �o���ʹP���#���������zt��뷈�x�A��L���vjL��"^a���a������ZPG%��������b���u%T��z�����4Sm���ӍX䂸�/.u�,�o����V�D���87�֝ }/�W�N��S>:� �g�.8��zv9hy�	\W��6����]s8�B���T;��Zk�巬1r�B�z���*E9�{F��?���!Ѵ� q�� �Au�5�.LG��^��.�_Ϥ�.r@�`��SG��U���`N3�3Vk�"Ԍ���f��0e\V	�|t����u�,>��[T��E��] �8��-�ɺl{����9���O��)�OL�C�����-Jɒ��XwQ;("�+jl�0�4�=�o��lB��Q���W�R�M&�hȽisn��J�]��"!��m�Jd`>󻫩FXh0�yτ�J����!��5Jy��S�h1�Pp�0�����/��N�|-�;�l���9Tb���:�9,r���:V���*O���֥R6
#��D�&���^���H��Y?E�5� �#_4ׁ)\�"�8��1⨄�H>�1j���!�#,�TW̆ �'P	�aΈN#�*9��S��[�	Uq���+��o@�׺;Ԥ�@����a6��"=�j�:����e-����~�/�~�sb���9/�
�����羕��Cz>A���x_^
M�T�1�HS5g cFU���NX8M\�F������50�^�Ѥ�@#&�_H�|o(��L��pԧ�q{���IA��L=��%*M*�t�B���W��+�[&�c�'/`B�;���m657��qd)�-1n�4�U��v�"P@T��/�����C����y�-�r��(|���d9B+�L�Ns��q��_9�aՌLk�w���<���Hμ�gW�I�!��W�O���{�����&�'��� p��B�2y�/�
��u҈ڞ���ӞD�򉋟7&lC�xa=���m�4��މޣ�oO��8�2����s(�5bK*k���#���f5|�%2����k����S�l[��W#wz���խ��B��r�[��GX�zo�(���A�f��a�}���[���h}��&�wF[޴6�M4�hW�p���y�������i��`X������u֦/�왂�M1$�M���H��n'u}
T,���B����~�Z��]�t?�㈓kNa�/~#�P�����E/�L���Cq����A��<�mF��̠��q���S�#]�x�wW`�v����"~����DX�dr���<�����Ȝ7�Q��S[�?�3Q�L�o_���_��*�?=U�w�bb�!@-��g}��1�}BmL�FS����f(,ي���FD�E�5L&I��A�G#�U7x��_���Z� pI��.Z�����C���2cfo>��
�X�}�����8ô	���
~�%f45��t���Y^Y�nQ�Q96rWD )��2�e����W<���_�p�DW�^���vB�D~��.���Wn_w��qZ��"~�c�y��4��
ea~$?m*��S1բ�j'��m�V�f�1S�?�(�rGا��A�L�C�.<��V��0�h��~:��I����@w�8��?/n.�M{���7�uwB1�-_�D��A�Ȯ� !V�#s�� ��y�����G@��j��l�7���ĮO�`�9P.��MGUi�����t:��ǃ��ub'Fn\�fvߔ���~G0���1Χ���g�v�8�UEb齟{��d?���]����g�A��Q����CM㝗�Ўqן
��$�9"�x�zfte��u�r��������*Т>�Ny�Q1%��<��%2�����$�m�Ʌ]���r��_v( #�EF����+d�;!*�׀`�.� \�2=�t���0�6�L�ŵ���M�?�}(�dAhE������͇cM@ngY�Eh́��)�b_�x�2��V/+��w�9E��ܐ_���3JuћW���d�$����p�y����MՍ����2f[l"t�BP{�j��%��j5;�z��g[.j�za0�~��2��\<�JCmH)l̨mz3П�z�v��S�_F;%Y�*;��& ��@u�=�m|����z���@FwkEU�W`f�&��.Q���WW|޽��j��K��c�]7U��t���K+�`6�"�9[�C��z��k0��6���7GLT�͐�-�8S��'N�[]��.Z�(�z����T+2���?��}I�!��3�S�Ɏ���C��hJA����7��c�4WM��M ����s7����E�k�㦅�Ӌ����Seq��-c�`2)���K��P
b�G��s��{�)S79by�+f�{�D=�KK�R�p�dkK���ua�Y�gWIk,�dt�j�|�&��$�©(�Q��9
tr��?�>�Jӌ%�`Ɇ�%.6�e�.mTF&XU� ���%�ʫ&o���3.:���9-�*���*|g�
I�g�#������SU�zhA&��@V/7mh+>�P��ܮ
�e��]ڹ��[��d�Lq˔5�OEN�fQXlxVHYEB    fa00     5d0��r��k�~P�����i9m-<F��y=��ɐ�mx.��/��FM�F�p}�:s���ܘ�^&:h�� w߳�D�������O��0]����Α�k�1�SBa�5��^�k�fy����x�K�M�<�<�ji���8���7��MBH�g���
�h����Y@\hI�s�,d"��1	�%�"Us��DyeSgD�.�,�O��@�K�C��F�G�z\���g��n��%Gw�y�粹� �"��r�+��$'lژ\U����D�V��lWW��$tŋ�xL��"M�4��va����ůMe��2���M+V����`Q���@��w�Z����U��~�_e�u�t�u(;˒2G��D�(o�b���{��P6������H�K`��ěa�ts�^}���+�å���sV�ͮ��tv�iKX����o=���!� b��a{2���'M�v�1�#�sH=��8���k�&+Pa	Ul�qI�7�]2�FE@��-u�2e�Gl=}�������F6�ښ�y��c#���?�6H�	��X�An��/�8V�M�O��悯��V~�5�@���&mn@�3�V�������1~�h0T��"���7��f��ki|��2-U�����QnN�tcsy���h��m~���:OK�\�mbe�$����T�*��g��Iz�Nm#�U��V6@��Nit��8�!Q�q!_*���������,�o�h��Q^�����i���[�o��)�l��Ō���ζI:ȻJ���D�4,�vG��>�5����a�xz����A�.@��4�<_1RW��_Zӌj��ٟR�m�
�������6z�)�s�i	���)j��f=:��ݛ�M�E���Go�����`Y���tq�����殟�t\J•��`JGs߼�1���Y���`)�#�E)vQ�9u�Z꛿	��f��r�X���òj+ �y��2��Ռ1��?1*C���?1C³,	�j��]�+�/�1@/�����W�;Qbey&4��5 �p	qo��w����U�.��a��W��g��|����-�k�il�0?н+���a�ȇ'Rm*��H�>�M�����V:-jMR���q�|[<qa](����u]�?e��f�a�4���%���皰��s��g�ֿ�J)���,�D��;���괜AI+�W�e+;�Ȩ�����=���!�5���p�V����!m0v���i�~_\�0��W��5��`aCZ:6-����e��7)���'8���|[u`6aK��J�ی/�-��"��u���:R�=m=a�aGJ/�& �M��xlV]�'��kV�I�5l��6��6ui�1��땬��r�8��6���j�Z�]��i�xV��Ϩkۗ�/7�QJ�����:���fv.>&v2�j��'(���=v��w�0����ӕ�爋I�\]��R�$RA#��U	}�������FޫXlxVHYEB    fa00     640TڝM����;��SU��_oq��4"�y�4p�4ᬁ�dX����hU��:��'���Fj�o\��JCGͅ�&-ȳ�x@1�<ٳ���Or���8��,"�o��M	x��Am�rz�,.�B,9�'C5Ս��,���b����KI�ð`#gT��7�IGt��[S���H�饒k�8����M�[<`?8��ިHJ�F�eY1��E�����w�u}�^g�ː��&[�]] q6u�c!�-�Eخ� σ�]e��t�C�:�L �c��V7P%���m{Z����SD��tn��F8b/��4�F�.�k
i$�(<��V��f@�]R�%بr�U�Ƀ-a�]��y-J��&�@�Gd�B��ʹ��V���h�3Wp'�krAf7e5�>i��͍U�ga�X����nFH�}�gS����fC��d(xM���{_�1+ 84��%��Z�����ޣ_;��E��l���KsTוyG/4�k��+³�%H�3o��t�	x�ّ���'3fm �omg����jܯD�)�a���J��l�O�V��V�H:�&I@e��5�R��tNp�q��Sk4���+FU>�]r����t�29�ƍ�}4�����B̠�gt��_S_E���4���`�լ<Gl����F(�2�F.I'+�m���+�;S���QE��y3&rx�:��d�����l��*�4��Y:��z.��^�w����L�.]�2S;��1v�PSu��-��6K'���3�g\	� �L-��?r\ɫdPq��e��� G)��eA��K.s����-�#n-��[�=���N�47��_|x*�u�w9��$��?���P��b3b<���)n�Nӏ�9(r"Lc|@�nj����D��TG�VZ&;���0j���6��D���.���1��e����7�.����Z��T"qjycK>ڝ�G �d �b��^!�.Y]��9т�+	�B�
�Q�V�
����V��b�P�j�����kҳ������#�#L��5�r��W*�bX�7�P�y�,���s>nq�=�3ߐ��e��#�&��� �[�~����"�21��P���MP�#�H�����D��s[[�g±�&'�u��s�t9�R� ���[���}Ԁ�>`��h�y��e�w��hW <양9H��I��uLL.�C�<�ET�.\��,	)g.����I�z�b�$���v��v��]KQ��0�W��z,�Q�	��u�HO��p��@J����t��7QE����|�'��M���Sכ��}�ΌE}�%��y\�AM�M�_����}�'�H��GS9�����;4 ����qk~��Y�u�~�>����#n���_ɩ�8�V.E&M���G#Ϯ���7�8`oS�"x����h�/[���E�����@C����Y6	O1Ί��ʯG�'�	�=߮)��b��K��T٠�3w��dםU�*����,��n7����ҹ8�����{���<��$2�3��	/t&��ב�t1����b�Η�[}���\DO��=�r!����ލ^f�o&���0܌4@�6�
XlxVHYEB    fa00     5c0dEȰ	�*F��`��,Q�!�^ctf�� �g�ZMmMӈzMV�&"��%wu��$�e>��,r:Y(�k��ȢFM�3	�0I�7�3�+r�~���	��#��d�[�-��$�!Yfᘊ}����
���I?B��>�JWԑ��,_�v�\&����A5Fzj�E[�|��������r�����4�{v����O[��IiN�^G@�DM�Tpt���E�@��ͽԂH�N���O�_��s[�z��2X�U��4=����x`�!�X��c��#u"��j,7xdv�!�����ጉ����J�O}H��@G�%ت�|%��?�2������"��z8\]y�7�0ڬ'�h-�I���\�F����hBG���%�6c�O�����罥�fo��Ճ,�f�V�Pt
e�^捶f8$�+��ad"{���N�a#ٙ����ީ
�1a�o������2��^�^�ߴ�=�q� �&���*��@/ܮİ햝_�2a����f�dL�*SIk���J�yo������wx�X8�����Awb�����-_���[�J=�r�����'��*b�A�I4��+�p�$`[�B��y���XT��L��p1/~0l��OW8^}X}�'�������`t.�Yz�A5')�>D�j���5E����gm����k�}��@J�J��O�Z���]8 ���
ˍ����A���m��`�w��Z��p�t� �����F�	�[��Q�koy�������B��f�9�7-N''j�KuW�ڦ��~|��z�̣��h&�c/!�&�v4���{�¤�i�
u�/pI��E�G�ԍa;��>�~5�XZš�夬G=�u����iY[&�
�&�|*�H��$�����ԓ��h	v��#Ybrǐ"fEdH͔v��`�^�6n�һ�3��)I��ţf���R�V���cm�'��_���Ƴ'.��ج��qj�y���$��$�4+�E�|��]6B��9W!bl]�d�4i99/�H\�s{.�5T� �{����6�0N���,�cs�W-���f`֖��k��#3C��+�J�'.�a���d=�iq3�,�:p��b__ÃF�ڋE�\�1��̷_���|^r��:~V�hˋ3�W+sg;�:�M����E
�`��m4þ{IY���6�APhJJ��V�9̖�p [h6b��
_�K�~2��GOe��a���>��j�<��0�r�Ф;f�H˥9=��JxKf@wn�����_� �?]�	���}Q���:�[u@E��H�od٩߬�D@������h`��2qW��<�8��}�!�3����@�;D�l�J��їo������}ѫ����HEc\�v��W�S�����
��VJ_��c��D��?� N a�L�Y������UF����PWK,ћ2��Ө���e���X�'���Bk1�ob�._�XlxVHYEB    d347     a90ImY��R��aq���zE�Y����ͪ ³�hF�S�m:�]�-0I��1��g"E3��Ŏ�i%^_!X
IY#�Q$@���<!���w5o����ڋj��B��Bf�z-ؚk�b&�������Q�����$w�84�7�"���j��'����lC�TH�����I�] >i��d<X��
����G�K��`B�%t~$m��t36�/�A�씟ԙ\˼�n� ���g�ǉ�-�����_����Ç����T&�X��ǚ�:��������{�%
xN�>u?���r�����i~^��y�Uɇ��.��HwMS��<|�U,�T��!}�ʵTY���xΝi�͛H�W��^����5cV�@�ѤǇo2a`�ا/x����)+�5*N҃�@�k^+/�m&���EP:�+U�����\�&�L��[�=v�9�n��$�I�߮3.k%pP* .Q�\4��s�.��p�x�;���]�g2��\0�=�"�3�C��~J�{nE���9>�|)�ꅡk�#]&4�#�\S�6aZ�a����7ozel�>��8I�j�Y���=O, W%�Ο-e�������4�wi&��ya��̒��Se!��� 3���l9���ep;��/�Ii�+�4(�q�{��S��B����p��Yk��N�-Z�q+%��C#'�����e0�O-��@g~q��
7�]�iGaq�J~�G#Ò{w�>pRl���ݎv���g�r���YR�kfs>V]Dmd��ß%��n���i.�x���%�o��v�Ľ�7Hi\�k�3ud���I4��?5R~ ⚖�>�w���J�����}k��p�	u�I�{&���M$�X��8�&,9���9A4eՎ:�.�t�hLh33��,����ǡC�����;(����R�E�1��<cF0VB_>��n�9��(^Эw�) �»f�h�԰��@쉈R�qn'�S���
.����(<o�?��X��?�)���GN�TZV�Tʶ��-��B���^C����B<��6��g�b�⵲ �F�Ȏ�p ��(*�@+� 2��͗&�Xէ�^*���|cR�hF�`<�L��+��l�~��Y�F�����b9�폙�a�D&���q����Ż9뙳�*2y~�-hVhy�����,�a���>��C}(�x�j����Q����sNDu������³_� bg��O�D��,[o��!Ǹ���G����|(��}7��V��\�U���ۗ�%�I��l���1����o�/�E?���e�t��AWB��k��=@4�P�~ʎ�	8ĬY�\4�?�z.���5�[:�C}���	�@�,MG9�%�Մ��4Č��_AEP�.I��������	��G��c�c(��R-�jj"�� QC�����*����D��"�3��n�Td�B��Rڥ���g�<�p:���;À�`{�[�!�P�4��T�}��<ӕ]�< �'��7k�������Mz�p ��.�A10�g������ᘘV,��^�I�'�U@G����-���z"���3y�qTv���x|+Gc�S�F���r�
�G*����w��� J�σVرڶ0�>p�2��XuP�n���}G�
��/Ҿ	*'�7:������K��.��,W;P����9V,R�a1����+��&1Ge��CCC��Y��Y������X�~��S�8�y��gj�R7A��U�j��f��c��媩~�2��V��ڶ[���9��`^�������-̕G@��� ����5��	�0�W�ŐI7.���n���5BDY��+�	�0�4��ʘa����}�T���
y�2M����u�	�)�U0i�>a�>�>t�~�Ȧ��̙� �V0S�:�͆����[[���q��B�e�,�r}=��B��[Sm��n�=L�2��p���^��7��TJ���nE`�.�$};����	j��&p~;�FQ^Elr��CFVIo��&�7ܲ'�)z�%:.�?X c`rxU�ܖ잋��!)ᑭ���	S�/���? �Mb�@j]�Sw��z�5A���!�o�H�ż�B��2v<��0b�/��`�R��G	W+��_��`���u������B���p�f��������w��U�B��%�;�۽g@����Ш�)��9�@!�\��A�
�⣽�c��D*{��Y<$���7�E��/���ɯ��i�o%^���6�����*�����=_��aɺ�)'�(|�� �,�6v�lj��HRx#�fv���ߊ`�LhC��M>��WP/�>�D�"n����H��	:�*�i���K���1h���Li�D�����,Iw�F!�����ӚφaV^ ���ф��O$'�/�/����.���;U�Z�҆���s�ುɴ�*�g�$V�W�{�� ��ްh��O^[v�����x�pU�������l�h3�n�Z�O`��p�[�[�(P�
H(�G @X�R\��ό�����lWC=9�9�� 
̿b��B1���E��W˪^�4Խ��9�-�)���
/�7���1[��9A"�¼��u+�Z�;�v-/�_p���N�*SQs�O���� 8��"gd�y��r���!��0J�4�E��K=�a�פ�U��m���>��ڻP?c�V�>'��nq;�d���-~�6�*�W�c��