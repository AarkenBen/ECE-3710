XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v��At��؂Ր�
�bt6���^ZIc�,�r�k��>|����x��E"�v���b�;W�)��p���x���+�ߔƢ=��8�Xj��_̞��>�Y��Ӕ Fs���Hu��G�LU�u�0=�K���$Ͽ�c����͈=���9�a����b�^�ji��#|n�=רܡ(��=�����T^�s�l�<J䎎iyo�@H�t$n{� 0�S�n0���Ǽ4�6��9Hif�_2�������mU4�t�p3��^ܾ�Jn������f�����&Q�q�l�jT��_(꼰��pmO`�7�����	�PUq�,H�F,�t�mZH�ⰺ�Y����|���.���}�>�.��K�?��Cw���tj�H��}X���a9fP!���/1�x�8x[FaY�����ιN�2Y�4^&E��b�4:8+d�j�x*�9�Tw
���GO��,!�q�������@0�>l\5C���$H}P�e��	яJ�a�x�h��m�&I��JHD����G�<��{�hܣ׎V�q�s�)��S�W�h���w�;��є*�D	;��3%��f���󆃣YO%#y�kk�X���X81,��Y�j?A\�����#+�
����T�;S��7"�r2�S��k)�S����k�`?�֕�s���3�QǑ�ŀ�s���z�}b���4��9����%Jl�ܦH�~��Z�k��ۧ"Q����0��b�P4��[�H��/�#�І�'j�T�ܟ�U�+ၠ��jjNTXlxVHYEB    fa00    1950�y/9���4���P3��������N�P� �0�-%c	�h���c�bRͻ�|��y�,�[���jG�����f��I&+-i���u�8Պ�ImB+"�Bn��[@�E��DrBm��I�U�U ��.ۻˬn�I�1��?�f�&�v��d�]�@'�T̕�R�~&ɬ/G@::�T_I�\���+�����V+�I-�@��j��xV��Ye�I�+�w�4��h�l邟��c�΂��i��1��ڒMC��2���bO=IXcI`�f�@�^����۾ ���L�#�#�#����(�5d�T��77=-��9�Js�8"�Z,����pl��{��"��B����u�j<t/0�x������i���gO���[�}D�z0�v��35��H�T��Mf��u1����8=��[Fq5�f�V�d�dn{]MFN���\њ(�/l�C�K���t��t�ҏaR
\*aZ����ZH�g�/�q��],z�s
&A�m'��(���ͳ�-����ީ(l/>����8�Ϧ
0�пN��Ɩ�ӡ�.�yر����C=d���v�-VD"W��/H�=��+N�MR��Ӎ�����n������tq�ǿ]i��n+��HR�u)N�Si.ز��>/��$�
��#���2��S0@��0?�'��|�ȝ���k����w�ž�P�0N�*�<�{�/9S��f�z�xo�s��zh@J��@_︤�R3�(���B9dR1�Zp{1�����.;�¶�,�j�P�D@�L[�(Yp�ݻ'kU&ˌ��¾����?������B����L�XixNi�8CP'�T�&՗�Shx�F��1L�+���#��k�p�{��ё���/�~��"��`��zn;f�&�XSG��`qJqu/������َ�MD�S}��Į��H�<;Ȁ[a��7`SV)���9��1t�?� ��۰ː�ӈ%�A!��R.�=C�����e���z�X�	�Q��w�7�%�i~���2��>����`Kd��a�+s/m7'.qI��h�<!2[����n?�j�<&aѶpm�ihW�4jh��PTwy'�z��LyHlle�bP% �.��=�}��(�Dh�B��G�DR�ylM�&��q{�x�4�gTڜ��V�m���0�W����*�dI���]4�D��G�t�o|q�^Q���%̱���� `t�
V�oLx��A�
O�z�͍P\%��'L�kD�,dk��FUPC���g#��*����s:�O��t���sh�&�E�vȲ�<(�T��=�e�Ч7�b�2	q�Q\�D�*��8_��%����k8yYNV^�8Nc���
k��-z������hU�]��u��{Y�[N�"֎�����R0C�=38����s�1�/h'5Y�k��՝пk�*iQbO�Ѵ��H)R�{\��a��h?H��I7�!���G}T��V#���P��� ��4_�Ds����IR�S> s[�f��`��BT$U*u���'���)roB2�s����E&ı�xNM�|9U&-h��[��9Y��yB~�MUTirS������Q��2�W��<��WtC�M����=�������Q1��Y��
H��m��[^&��T��3L�c՘Ҵ��~�n���c�ޮ"Ir�޴�8K���'V�`�P�ēQVzȧ�+��_�N$F��ô���1҄��ݵ@6:_"z}oK=��v���?lWϐ
�g�'���\��n�Q�~�>5M��'s��<�IG&'s�ٻ�]Y�ާ�r�oǸ������a��RP�O�x����d-�U�@�@��U�>?�.��*U�}�~_�;���į���VOt���TT�@�G2o9�2��������3�\<�wJ;i���@f�8;a�` �P3�beg����=ˤ��\7"��_@t#�v��g�O�D��Gg���}מ�n��gΖkvq��@�Mg<ؾo���̢�&��m̬''���\&jx5g�#8��!�0P�&w)�9��H=�A�
	���,���7�A
�z���k&n����1F�H�NoXU^Ƀ0����h �6`���3�TZH�s�u06N�`��f�\�y��S�h��md��ё�s�ڰ˸8v\��_����;�z�`��Y�B�c��K��g	r~%�@�m��Z�?j��Y���	&�f��p�M�4R�������bp��Ϛ���g��Hh��>�Fɍ���5��r T�fzpx��P��|V"�?�� ��1༮��%����=@1~Є������$Y�����G���XcӮ�7��Cێ@(-u�RGB5�rN��ţ�%�t�/���O�ȃ$���b]�֜\rB�{��3f8�9���ư-�2̪҃�����v�K�.���vl����.��$Fg�0�|]�S�ݵk}�����Ld��~��y%��s�yF�5Y���$b�H>t����%Y,¢o�Ȳ�]��S�~mQ�J	�xVкKux/��J�U΋R���u������v� �����SQ�������_����G���4cj^�N�\:-E����]J��Ň6�4R<3u�	��gИ"�����d#�a6�-㮷��'ʘ�5>z��.,�g��29�S�	�jq6PϹ��,R�����R�pz����-�Y�n�����uE�ϝ�� �_6�GB(��q~���@�R�X���ߖ����xq(��J���
��T�-�̸�53�F�����1�ػo����(��
:7�XD�(eP"�<$nn=��U��*���҄}���38bQ+�S2�q��BW* ~T�@{����Y��d/|?Cw�smS:���\J���B*{���m��_��;#�������9�O&���m��T##{Hy�a)7����M���vdnQ�ӡ�7��!�6���hڰ���%җճ��j���,�[�����e��^���Ҭً���4�b���T��N��|kA���h78��>fa[��%#,gg�n�>���˱E'��F�>Z6f�!�-�"H���K{���|��ld �B�Ye�,��uJX�4��_�ʗ�uQU�U_�'��O��IC�������"�X�J{���W��k{#g_�"b�v�	m3�}�˝�RE1R�����+7��3�O��=�[���Em���ch��r���e�[S	�:��];�!�6�zZ�*s����;����ӊbor��
�����2Ŵ�3,;���+8 �`wp��NϾ׀�ƅ��g�â��W�뷟�]��	S��՜��Ckkz�����x`�[_i}[�sB��v,3�_����e��7M��P>����j7wwO�7V�!vL�hU-�.��L90M���w������N*ސˇ�39�k:[������Ӏƙ��
zp���^��յ,�\�C��߶�[^��C����C�sl*+���^����O�`��M�+SJ��d��C�6"1q��x)��W���@h�`���Fqjn��{ `P�N�~%��D��7��!��شMh$ލӤ����RH\��D�0�x+ܬb��>e�Љ({��j�)�X� �B�t �}�5���O+��kpl�1,Q����V�7zQ��.#{¢{:dӒ����fj/@~=~n��Ya��G�1�=��������RAªC3cIeE%s@h�����;
 C$$v㣡̇K� ��~�t�&�^2�BЭLx���%��Pݿ� cd��3�+!��к�����c�'3�6JG� �L�����S�{��Z�)K+z���ѥoX�a�
氓}ߠƏ����T�ﶁ�d�c뀽�E՜w� #�Zf��*8�\�1v�`��K��|���h�*fK�$��@��S�Zvc�&��hJ0��`��1n��4(������|��uP�6����b��bx���[�!T��Ƃ�XK�+(�Pڍ����/	GE,b��w�F�#WI�<I�[ҍ�S�ߥ�NQ��=^ҙa�<��X�xm��pL�����Yr�4���]�=��ǡ
݃
sz�U�z�uMpB!�Ҭ��wo�|"%qR3��'��RC"��I��Ԍ�6"�y��=���%.��uf���P����R�W��!��p���GjX�+Ot�����'�h�.~�M����*V����eToF�g�*���K@���y!
K , 
�Q��j�A�0E~,�ÂU񝷞�0q�N7���jR&�j(�	�\RU�lR"�@�U�M$����S������S_(���/�-�� �IM7���3\��vb�9_,�fr�GS�@���<�ω�ϒ����<�H:r���>ՠڛts~+�r$ S�=;�e�W�,�Wc�(M.�à"{��R���ו!����ˣ)�/%���Hg��,�0������Rba��$��n	ӱ
b1�v�ԣx��9I	��L��$g�w��Y˳��G�YZ%�̘*��`�V�J�zHs��
,ƛ?#�hD�.LX�p�#h�k��}�����dfd-���b�����J������+�)in�'�n����a�>h�ɋ.�q�Y>���"��>�$M���E�&jL�3�_��������d�b�y"�,�VWY
f"�襝�F�t�J�l6�ڽ�cBEm��&c�$akr��yY��kɔ��B7y{Bز�l���\-4��ڤ�j1���D�@3�uO�7c�y9ۿ�PDg�]ك�+=T%�x6&gy, ����#��B�Vx�4������?��tO�K��/��������ړ�p�4f�~��g�d��[��q?��Fg���'����a�w������i������eO�Ⱦ�LC���tS��藆���D�'�hݠ\j �ͺ�IK(�\���~t�. F�Jy��3\�Y*�Q�aD�ۚ&���W� ���fih���Ԗ�O�@-�uDv�O�0���?�@v�IP�Z7�n�' ��M(T0�$�����$���1�W��[KK����L�JZ9���-�Zʜ@f�Gr��f�2B�>M�x�;I/�f��'��E��7��.Y��@���
�0���Ib���GQ��v��ņ�Cfm��α�0fˊ� H<$�U�z�ʽ[��X��I~�U�wso�[j��i��N/^a�Bv�S���X�#�Z��<��#-��Z���)je�~��7v4B4�~�DW���ݥ�i�l``٧8*RN6�ӯ�{��o�f���S� ���

��S>BZ�Y6q�A�h �i?�?��cY5ʟ�z����'�N�y:�8�8o��@r�T�����[7ǿ�S�Eol��=f�y;1&Oϩ�x
��#��7�;+v�oV�z�IM�H�	UY�Z��jb��SA7���|
(� m�IQ֤�0�`��.���y��9vv=ң�&+���]Q�Ň���dSj��@�ɄR��{�[�c��O�.�S���E�y*�.��Tnb�1p�T~�c��=�<�G`q]��� �C /����[�iT�ժ�:P���)�ڌ�$���}� �;�n��.�q���'���SGi!ƚ�~X4N;�$�B���C	��)D$���^,��K����9ZV��D�{lfn�ef������j0|%&q�;Y�f�u6�}���9P,�$�1����z�
��`�"��
F�E�0B����D��d��4kJ[x��~��%�^LMZ����E{�"����-1iᎠё�Ǳ�]��A�K��A���se#7�.�ዥ�R�ۜbz�A�Y��Y��ٖ�
$,#J��yՄY�hx�&�S��x?�,"L?QD��:n�/��m��;Ma�}ٍ�:�|����?��M��	�Ʈ�{����J2�KB�}T�+��f٢��<�)�)�a`�t5��1I��gkm�n���|��O���=�r����N�����n�
1ߗ�����g��
��G�Z�}X�.��w�ֻegw��Y�j4���W�f�"�J�w�3�tw�!��$`9]��̛���i!i_m� �-�e��X75��vXH�8���7�Z~Y+����PB��G��܇�F���{�Z,?�VrB)��<�j�(-�Ц�":���[ ��y �o@��,���i>�(�p�*5ߛir	J�r�?��:��x2���0�W5�n����@<՛�ˇ�zET
����r�D�[��]b��M���mBP��"�Y������_�=�f�Bt�ELZD�	5u9Eb)�����������d���~�!���x�R��ď��,��]���OT7-3��[Q|�۬x�lrXB�K1�&�jƷ�ܳ� �SL��HV�xʥ�|c"��L��\��X=�?���<7�R�9JM�\O��97�:��t���P������I%lh����K��bf��=XlxVHYEB    fa00     700(N|~�Y�.1�-]WV�X3�4����� "�H���vE(�E�l��=8�����3�׎��:m�v��vt7i���8�C�� ��?	zΛ�Yg�d��@#��"����	�9�4�#��
,R�N��� }�ﵞ��.^20I��Eu�?h��Q�O��s޺�C��4$���N���̣�l]�(��{�g�l0#Z�~:�XVFW��U%�˹X�8:�I3�^H�IX�c'�4cXD ���x�/���^��g������"����ݹ�@5��4�+�e$��Å����hZ~_c��'e>�Q�D�@��'�	���`�)(8�0b�5�g�/���f�hb��sb�u3����[wz:�A8����Ϋ��K��vS�k��X������L?�`^�>A2R`'�[����V�BJf,<Κ�)@�i]0�t�a��D��mҊ���4�z��*l��z����nB�������D4����S�\ڣ�a�̇�
%8 ��\�*y���?�~�2p�J�߭��&����HY1�ds��^��D����׿��;Na\聢��!8l����;���s�@�iŲ�Zթ��Wc���6^x*N@ع�a�9�ߋq��A�'ز2^�A"��d� �X���rx�A���|����8�߅�Au��ی����Я�s��?�
cS�R\Ј{�¬���<�G�]��5���W�r�1�Cp� ���i�<�y&>r� g�ΑC��vPn���0h��>�O^ ��NܥQ���˥�Bl=_����kwc��ya|�_��t#P-�"���$ hD��X�߯t�aI�?Ɠ���լ�qk���sB¸�7ׅ�0I���ǧ�֟��;Uy?� tڙ����3n���B'&X6���d
gq8�X�Յ����8���:a��`Es*��+ߟb�f_�ɐH��V��ҁa�=��@�h��ЉIN�O��!��p0��O0�=1�v��z�d�;�؎-�:Ϲ�m7�(Z��^B��oB_H1?!eE����7)p}��`��3�1�Gճ%���������\��w^{���7���j�k�l��LM����,�]�M����B�leYk���RT�y��6���@��S� ~�F4�ǌ%3�]��
��˶�)#�}cz�x7���g86� 1���v:{����[l���BIw�|zT˦\@���M��c�j�ȑچ���뭕�VSk��3�E���Wi�[(��`�|���r<��Ws�T7�@�1�ꅦ��r��G�`����v���v�H�X%��K���>�pm�C��12�k���'���W"��Bu�J,@TFv����`��2D��cۑ��(��},0N�9�޵H�jDU��v�u����1��\�i։����>I�.����o�71~['�cb�|��x�!S�n�dh}A��&>��m��~%�.pAXw�^CxԚ� �A����G2���>�Eٻ)o>�~��u?����7w5�ԃu��"a�̷N�vz�%��,FBˠ��%˽������L�QF�N��^R��T�M���XH����EZ@MJ(A���G��Qj���X=*b����K���{	~�Ј�X/B��0_�ȯ�I�`��̰����񀋥��I�m��-I�p���M�S<�_jFQ/�`���ݍcۗ=���"���IA�s�.n��D�|�Ĩ��/.���a+tUT�˃W�M��2;)�'Sk07�rN���X�^�q�Hv㷮�M{7������z,.XlxVHYEB    77da     a60��&M��_v��zs��$S��[���&¸w9���l�� ���pl>yֽH.[`c���x�I��f��twk&I�*�{�;zB�Hw��x��J��ܿp�v�[�Ӻ��9gU�4׺�10�Oj��$�4��������@�]�s�N��v��[�+A:aZ>����xʾ���,��-��=�|I���g����8{` b�v�� @ՙ��|�b7�9�=�ɓ�<@E��bm$��6���oY8��(7NX�֕���(IH�Y{"8�b�='�!d�>f}Ǚx����@v�Ҙ�iic�i##�N��(�ǎ 1��τn:F� �Y���zA�����DO�bX�^xУ�L%���bA�oW�N�3"��1�}��u�"�yN�>J�-&�����~-��h����0�J�PO�����=D�ф�2ܿa.�ɐ��(��BaG����̪�#7�J_�1�k��V��k�P��LN�rS��C�l��O�\�/s#�ێj\��2m�U��ipq���#�w������\���+1q~<���ǀ,r��É�u�Z��Rи ��~;��k��?Է����5��"�Q}�J���0k[�) �#�:N�#i�W�[2�=�Ϫ�t�:&��@�4_O$�B�d_P�B}_�y�JWx��}��J@Sh8��0�����ޓ�J�pCm����jSf�+�^ڢ�П���3�]V�L�}�H��[���q��t��Q�\ �S��f��G�Zp�Ɗ��/ߡ�A�g�LNB@�,�	ay��B��,�-;���ݢN��������S��r)��i��88�Ɔ��`{@	P��ͺ�	���>s�O1f�R!o�K��2O*�!<�W�sU�� �C�M4�4J�Sē˨F�=�GC�i�J��������I'��Ɍl��T}j��<K=���?~E)�E	��w�G̑چ�*R���4����>��;Դ^�wSd�7^YtU��*�Yuݩ���e虂��)� ?�p_�xjB�]9��,��1\�R;E)}P>�y��5�Oq����ѭ�~=*�S�7��qw��]�谒���;�����K�N�4��=Y���p�h�FA��'>��C}��v���;�0���	�.:�0&�!qYԘ��f_&x{4+�B�$̼~a���]�hQy$O8=�)̠.W�S�-DoԘ�� m:k�ư�k$�0�r���p������3z0~p�":�mزd�/u�`�E)�N����3Z����?�C;��9G*�ˍ_b��Q��p w���0�5�M'�����VqX �"���cT��55<jU�ƞZF"j<�|y���)����a�ڰ���W�,U[	>>IR'�@�Lq����C�4���q	��NDԉt]���dd�5�ׁ�Y�Ygq-�<%�B���w<�f=��Ҭ;5�,>��S��ӈ����w������B�r2�<�����E��C	+�&�G|��?*`cʿ˕Y��I�����X��X΁-�$0��ި'�)F�Q.P|��u�cy�-�$�W���N�#�7G���t S+�����8cZw��4����"�T����G5t�1GYcs�Vӄϫ�����zв�?��l��a"%W�Цӵ���mFx�� �8�2W�}�ֹ�3�f�@uea*I�j���K1[��Ϭ���ld�����`��^V��&�s�?�ݎT�sL���	��*�"k�5=���!�ݨ��!���C˱2��w�>N��,�fNV�^~�w3�~K�<��.�?Q������]䮛��B����N��6�^���K�)3=��鯂`��&U��4%]�S�k��L�c\�V��p��7��bz���;/�Ԇ�_1���{������ئkVrG��q��'�V�J���X6�fq@'x�[�����Y���3MX�T��`��������0���ܺ,Stvu=��a�9ʮZ�����x�D	֔�Z�Ϡ�R�bHF�	�x�<�� �y�,�"F�߫�� s�W�����:/�t��Wl)J%�A,:�/����C*Ԝ��-_�ut����.<�/[;f\�GT��9?
v]�������a~3>����^������")Y~賔8�(�$���l��3Mwo�c��D�Ǚ��v^�Qf�V5�)N+K~�_��w(F�^�UD�:.�!�n2S�u�Dqp�g~�_��W��9��!G|�UO�C��)?����3�V]��L�PX���$�b��7֕�h1�ؐȲ����'�,R��O�z1E���'����e>���K�4Kck�Rtm�?5�X#�����Z����?�A���2U(~���~,��n6I�y8�N3����w�x�Yq֣������ח�%$���4��ЖD:eD��QN���s��/����&G[��sV���}i�E�
{p��lU+Ɵ�.��$���2l�`�)�3��i���o���Q��zr���07�d����XO)�;XT��e����s_P���~]�e̋������^���5l��(��3yȽ��,�Ѥy�Yq �h�>o:�V�P�5G�;��a��ͻ�\��Z�b|� E���_�Ǣ����&��4L4��-VW1Z1�5�Uk�-+k�Z��]~Kv��fc��onȑ퇻