XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1���Ri��AEĤ!vy�Tލc��ʗ.L*�]�t:Ob�\��P���-���2�t�`��d�3��F���3��&�[ }&�TS�2�U��c뺯��3�k�ZWSo�C�OS;h8ms� a���h�w��E.M������<�D���#F��oA��'c�m�U� _�,'��vJ�����@�$��q<9��7��Z�vɻ�6έWSa8� M��Gf�����^��rߴ��dT]W�̖���6�k��R(�Q	�ˋ�5�Q&:�LZ�x�9�%��fd���
]9fx�Hj�F�f�_xd����
��i�����F����$��sn<-��u>R[�\���`����6��T�h��f:���U�L����q�i!�X(�37��v������܅�Zx��Y�|01�v�۹�j�_�_j���G���Osq$�n����u�u����_y0>�H���������1��;M�yyZ��ED,|�4�F�,� @�_��w�+�� ��ٸU�R�N�g�*�e[��隻"w��zi��qW|�!Ԑ<5r�o�F裭��]��O ׼�ˁ��Y��H�ة»�v����.$� ȗ���>9B�pĩ���k@FJ"Y+̘ �k�5�7a!� ͵���ձ��?�l�gW�u�;���@��C��&[a`�����K��ȍ��!Q�~���$e<�{"2�JݑNu��F�Ha���V��6m샅�$	șB�*={.�OY�M*����C16Q���*�?����c��*��̐��%UXlxVHYEB    fa00    2910`VA.�\�ۇԏ���w� ��ɇG&a8�@_럧����7�hMvT�6�w>�"��-�edp�a5tOJ�4�Ց_��CY�}vx�8�$�|�M^�9s9{�p1�!4i��D��p�%���hwa�HBD��*e|�q���q����lyHq�Q~���7�"�)3� ߴ�=[�ހÒЬ����5X9����QC�^sD������8�"��XF�6����g��&ɤ�̱
_���.w�3ݪk��'~rU,�1pH/	$�������-;2��<Q68���
i���,v=:t�������FfJ��<�{��,�5�(_ ����c��c�
�a<���T0�1���؂�g�O��̭!�l�LOc� o�����B�����=U�P�8HK�k������~մ��R�?r�p�$���%�ĕ���|�[��d�X�b9wl��.��}�7�3�Mt|T�F�T�Dy3�3d�@2;g���c&������:<�s;F������f��ý�J3�p�!P�E>y���h�Hb5\�~�� ���2�l7������po��ט*Ɲ���E��̻���Tb��g�~PV�o:7��)�U��䎃�l��_��T�X�+~U�|g�pd�R)�T�A�E�2��0,@o��֜�h������6H�	�L��+I��c���O�9��8"[�<�*���ذ���Y����u���+T�A�wc�M8���JpM �U����+�p�0���	��o0c��)�"ߣ� =8�"�y`~�ǝ��HG����z�� ����D�i�yn�����s<3&ҊE�T?��j�ڍ��jG>�^���=���H��?⯠�$]]�(@RS�$W�^gN��Z��kW��fg4F�`���EFe��4�Z��4�򌚬�K_��^^QY�_!�6J�-W3�[w�e�v�QV��S�����*c�:����Wත �7�
l<�b+��&K���J`MK|�A�Ou�75�G�i�|��w��h���ŖO��Kx����������Qהt���C,2\1�;��̢�X5�DSLVU�DxfFH�M=�y�hA��vޏCPNt%D�˷��U��Xy��{U�LD�#wi���/�Y(��Yw�܍���_oD����eL�x�Oȴ�ήO�}RˆAƞR^�Rvv#ϴUM���P+I��U�ow�~���|�H��?�����w�_�E��t��dM�&Hkͺ��������$������/{�S��$V�?֝�s0�l|�y_H_&5'VX�elo�Jz[���_�_�:H��S4��g��A�m\1�'��s��J*�r�D�3?�N��[)ɓ I~��	��V�>h�t�%}z��G//hD�Ne���F0>�7�r�����G$l<�K�{��P����J臵=��$���kk�1D�5�mȃ
z��a,.d�*aGo���w�����jǋl�s%xd2�|��?|M��waG��x��iN��_�*dUOw�zS���Dm��ii|Y�')���wa��覸7���˰���{sr�Ceڕ'�y�]_��&r2���f��t�G}@����㴄/��T7S�N��ź�q H`�nT��l��<wG�=j�'�+�@�~�8�7K�DhWAH�VYn�m�z$v�^�G�ZU���5n��CX��=�D�ƓH��%��'�^��/�>sv��jD�����>�T͛j˞_���bG��4�������N ����Yĕ�K����])��O��j����0Ha�����͌�K���%�5r�n="+��+WgƱJ88(Uz�מR�\�|��^� �Y0��F=q�q����Y#�_6O>���v�� �鷢W�NF'���[b�������&�B�8*� ��̘�3bYw�G%J�Ƶ"��g��S��p�\��9?P�&Ԏ�� �^��Bm�����O�W����*�I*]o@��oΧ�ޮ�j�-��5��h�S7`,��6I+,�CO���H~�(�� �5k`)���g�Jp��D�8}��o��?�y�ⓔ�PS,�� w�7C㥟*O�S�*K��qh
M�:ǀx��~^wm�Nq����,����"
����ݿ�y�%�"lc�?�u�#K�1�d�rj"�L����B `��,�Kb} l�TƖ�p�6�Z���e��Hi�_K��y7�m��2��G[}�MA9	��׿�� �L7�7+$0�������w!�a�#�f�<�\�r��_v��&v,(흄��Q�g��i����i�|\�
��O�6�n��d6^7���tm��Q^-R*�M��3d��$��M��x�%'�~ P����!I�|�Ζ�K��b�M��]�)	'����a��j�_�C�w'=<��+�w�$��
Svh
�1��\#xF������r��5��bz�����@�Y���3��#�G�mb^M�zxn�_��T�\��5a����h�g3E}�U���B���T�C���;��!��)V]��	��/t�n���#Cޢ�r�jQi��XW��M��(;�e+4�X!}�l��q�|��àΆ��-3�M��+>و���t�;�"zoǷl��z��ρ�)��\��C�?��"r*��	�5�½C�����u���rB`N\=g��Q���O9�$�/;*�$���!�z�P�)�S~�w.zC�;���tc��e�%��*�g�	�����$3�	���d�<S<4e�ɂ��&�Q�[�5ɢ�XSV,���mU���:�z���S"����:%W]���c�T�����w+�NJ7�Q�Դ/����
�? �-|jI}��W{W�{��r�NbUg�9���3?�^������c���lt�(�����' /��˦�� D_vܵ�.~՞�b)FeC!�̸ޱ`&�7�K9���h9�� t�w�/��BEr������ �L���(�y1y�&�3!����S�a�\5PT;�e����S_����H1&�=I��|0@�xVWmfL\<�@Ympe �!U/=��Q��0���s��r�����oD���O�xwP?.e��2�@�s�n��L��{k�����=�Z��Q�D=�L�}t��&F�)m�Y���
>�ږ-[�L3>�������3�F�z��D.$U��bc��k{%͔�E}4iI���Yj��v��T
��'G3!�Y֕��"n�����s��������T�v[ �HUd������\�`�F�L�TR ��W.GN���Nj~!=6m�o��`w���sۗl�l~�����r��0J�A�2�C��n#"�C��k�3����_�E6^9���)�?֪$P�饼ޓ��!�GǛ�bY��Bo��N��f#��h؃m��:�� ��;�O6�կMbx��¿n��rj�F9�`�X_dv��"�]y��\�|��p|��$����?�gk�� 0���D�D��ԙVE�b�k"y�'%��s����H�)�I��-�Νϳ�b8�{����m�s����uhڼ�k�Vk�3���P���j~Jr�
�W`�� �I��#!�'��e�<:E,�^r
�ᄳG|)�����W��j�z#�\ɲq�5�)Me��+r���޿=�:�2^v�"��/�V��:Pi�I*>�9ѕ7_y�CV�,bq���!������b�5UO��v�G4ڌ�0A4s㎛X;Dr�����d��7 ��ϟn�M��λ���R[���X�
5�[�M)�p�Dl�ۯ�Q�q�wM@HB��`ڿe(EcG�~�E�4tm�Z�=�ñ$����ǝ�=�%59���]�$��@D���ʹ͍ȧj� ��h�|�st�Y]���T��W(�P3UH�D2/��5�1��.玼�b`�K�x���9�L���� �����zD 
bx��{�7��5^E(O�i��2�-�ѯBVrL��)���i}m���j��|��,����l��&���JF����4}.���^�aQ��Y��V��+��:��>�ݚ�߯T����\������*����޹�<mB�C�@m%X���1�D�d�F}È�����o_ ������x"�~ϧs�@!�7��+���Ώ�=��N=u���<r�f���{��fv��xk�_c�
�J�$��r�Iy=!1����-�u��w���f9�N��w��-�~��2��r�� ���IO�3�T��9��T�����B㧔 ��\q��� �V-��u���C�Y��.���̲����4@�qA��Ɖd�IJ�t�(�dm�9$`��OFb���n?��D�>�A�c]`�(����.uA���i\ճW��"������~�i���؍�ί��N���>X���0%�'��6�}a�!mځ�zj�l|�!`�EۻW(Y��'q�^�
�����	��t��{M䂌EEy{ڶB��f	��,���s��V�NH���v��D�y$�㼐t�G=cd�sg�n Iԗ��=`�;��6t�C� B��q��a��SzI���*d�T��~B"��욒��E�� �I��S�C��%Dy_�'R�vH��۳?�ZH��v�
�<|���IN���sْ�-�;�����LPg5�Y��+�K�l�y4Bjh�u���t(U�������]ΠO����<���b�KU)���R+(|�Р����x�`��c�v�������4N�bX�uL�|��$P��:���a�_��xhJ;��Hhz<"y.pQ�R����+�q�Y�wm�K����u*q��;�lQ����i��h��2"��)����W�9pXCYg5NZ��b�	�0�)��H��,�f9�����b1o�s!�"�[��:�����Q��k]0�s�����a�n!��!�h枢�h���w;�s��c�	��$p�T����>ʬ�=���7L��Ŵ&�����'P�=�n��k�#ƜDE[Ϛ9�g���Ұ8���eM�qΝ�������2_��=�Dm )}�(ס��W���e0Q�v� �6W̃A�>�`_�N�P��é��*�	�ny8U�O0��Fk�}�4|�*!sBn_�Ǘh4E�V����`��/����=��֫��s���=��h���y�?����.�%ƭC�+�j𛿵�4�o���=]���S�<��2��2��r9g�!�����y������eܐ�U��'�*�5��)�Y
�9�)�m�_;�w����*.��?A��|!�����դ���Z�M��Wy��g����U�A\aŧ����J5���Znl�ݔ(��w�$�����x��gv�*Y�0���"2R@��ф����G%h� �� ���`����0[��$˙��������Mkxr|k?[�N��( �+ͷ}��>�:����!-�x�S+|֍�J�n� `/ԑ�}��;��X坩P��+��� ��/�BQ�(S������U�y�v���T}OX-��i�#�Ҏw���ğI,kz>v �<"$wl{��?�u]`�;��T��$m�I��W���Z���	��(Tf��xGʎYJӒ���T�� tV����P��9Nj�Z��Zmy�����`t�����h�7���]�blD�������z�`x���9z[�f�%n���'��/O@A��kJڹ��.Tϻ���3�A�g=��5]�r����d�<S~�q�x�do�nk�}&ِ��?Sa�ƑT��݋��">r��8j�����v�G���՘���@��s��/����$k�e�)���<�z~�����8��lT�h
|�fd�J��7�w�sv=/40ï�y�as��o)4.�R���������50��#���j+��!��K����y�&Y�ȥ��#@��UhM��eM+H�����>Y�ʟ� ���T��S�g�=\vs���Z�6H�C���T�,q���"(`�М�%IM#W��)J�S��P7�k��stR�j`�6�`��Ϣ���շ�=S��:�o����܀��c`T�a�zTHc����a�"��Z��Չ���.�4�tI�1܀�|�{�j����jm�L��Y�f�� C#�8�x^��O+�f��m�R�TM��pI+5�lʥ:��>�A�G]�vO�H\u�|�\�C�����.1����,���I���ݩ�\#��l��^��\��:���߀G�|*��ChQ����y����f����i�}��r��;q��"�bq�;�]�/T�l�ī5͖x�н�C�_�l�1�Gr�~�>���l��u�h~��2����ҀvT�O��AS����E��7ɇ��_����N5���[_^,�!���ت���$Q`�TQ�q�<���0L���k��ԙ�>e5TW��?�,�������㉙�-����� /$�Խ��|�r�eaRq!��fè�bC����ӳH.���'��WC��١f��`�!�|uy��5�P�����q1O�
h_��<�o �s�'W|��������I0k�Dh/���	Aγr�r����Ҍ��_������& �އvT�R�t�U�+�S�I��7�NO���zwb�k�%%>��X<z�eF&b�n��0%ܩ��k�*h��H}���ǩ�U�
)w�à�Y�`��wiJM3\��`p.�-�o;yrp�[�Qp3�^d�};��8�ڈ�R��J7�sf�w������oފ��P��Fp���D�Nڄz��z�	��=���ޙ��7��1������01����'��Hu<Cx|������@�M����(eWBw�I5^��j�:�-���Ԯ:��y����
�:~��F
z1�ѩ������~v2�%Rvw�UЇ	a�/��s�\�����K��0���0�*�cP��+s��kO�`�����2e_������a�R�h��ko��hm����^khP���mU��A!q�cB$��������S[u��Ш�#��`��l�pY��a(g�yH�^S!�i��;( �Q.ݠ���I�z���B�G$24o�f��e�,&��^T"Nop�;�\�r�Ʈ�@����^�	�F��Dv�(���; _�,�xr�llBF+��A~������ue�Z�N�>(}���s� ��d��� ��e"H�o� �Jy3��&^3r�9ӳ��k;�S�H�%���સ�mg�m�Y��^P��`1>�YB�us�蓆���a/'��1Qx�m��W�?5���!2"������lնN�ɦΦ�HR|���
 ]�!iP5�t�zb���hʑ�����\����޹N�G�tʹ���?��E����J������ ��A� �����{�D�0���x� |!G�V��t�.=��3���)�������,�?��K�q���ڍ���T�֐ț��ƪ���6}�U��<H1'qWHb0Q`dL454��y*�yถ�m�8��W'ǎD{qE�Yf3�2���-�[��o
��A�^m#3�:��G��%�4���|�w5�7�4��HI�@�g���,���I�L��BcC��V�a����g��qS6��r��ϭ�lP`��Ȗ�	<�領vQ�!�'�D��B�W����&���'�o|Ȥ?%��5�D�F�]fl���^In��h�<dW?�����n{�"�y\1cmV�������_�Qn���!���&�Vq�q1N���y���H�|����R7{��	�-�iU����Fu���b��3��2�ݛ"Hh%N����$��0j����7��? M ��<&����.��tC�	��CL|��v������3y�Ϙ�UHY6[��K{����-&�ݦ��P����Tۈa��|�-����3[��
\L!�5�[��ׂ�� J6,���{,<m7;Y�"�ܛL��$&��q����vN���\�5 �?��m�@����rlC�U��9T6�� 0{C7~SƷ��cO�f�R��	~R�q����F���#R$[��^\�i`�����ئ?H�"?��* �B/����D-gc�^{���\���t��A�	��z� a�ݨ9�HpW�@U��ܻ�B��Y0�R�^~
"E8"��b;�����7������O�__{{�ʏ-��_��@��a����D�ןy�B�:6w��ӏƼVS�/Mͪ�D7���}��t
9֗z�t��taP��B�e�# �x����y�1K{������Hu��ʅ�=����#=�3	]�K!E'�\�4�!��w�&�bI��;�%���L�C����~Yv0W�@G�|Z�W�2��
���~"Q��t�>��'%$E#�E����N��l�(
�7��N��a����E��^!��}��gpx�-��6th�����;�9�PT������w�:�ؕ�W��_��θ)���*~c����|�n�$>tFÒS���.zA��/xĖ�,�{sM�4�K�ޮ)�r��vW1�Ѳ�ᬔ|Q��&�8/Z���t!����E�:��J��bѕ܄D�~�{��6�j v�Z���H@�]��U#dݧ=�Z-�����o��5��֝�O�f6`���x�HQ ��q���<Ѵ�J�yQbY��K���L�KqU��j��	&8�6�>��x��H7"�T�"�(�;'���r��_�{�7>u��KWX����0;���M��K��艅�J{*�̕�L�QCY�m��A��z_lU�z�H��Z�(N���>­Z����#�hP�����}#���rw�,�A��5B{�t���;��cҍ4j�OgJ����\�~䏮f`$�Y�WZ�+��O����F܍�q��"*�XI�J�a���Ձ��} �n1��Y 9�嫭&���E1}��j�K����/������u;���l�x�Duϫ�$P�gb�!v�2]2�%��4�O�h�f�;T|E����x�T�ɋ�=�s$���dP8͒�$�������P��'P�8�t��_�I�����k����EZx3r�Wj��2��f�H،�,�	cV�^I��=-	�"y�{Z?�R.	*�\K�x/���:o}�k�Rp�7TɜE��%�+X��~vQH4}<�D���3>�\���y�y�j�M���m�x������
�y(�h�O��j��ݯļ?m�s��q�.��^�X ]Z�S�6-	d���(n#���f��P������i�H�tI���s�}�g��!��l'�e�[����o %�.
�>h��O~�������|_)̀8�H�dip`���B����V��̡#]6:�w��BvJ)d ����c!͑@/=��}����Ec��9��Z��D����l���Ա���R���}p{��V`�K�e7%��� ,	�����t�/�56~�>�N���!M�Q��:18����Ԏ������?��P�Oϒ9������#�v�%�m���`(M�k��He�AC�#�����Z+5��#�ea�\�?��ـ��7k�����7�';�g��{��$�	�>��xꆷ&$�����#�6��/���;:�O��o����-�cT��=D��MB;L������XeUd�L?E�V+�	d�|M1�WHP���{�$i�V����BE��`��f�F&�C!��h�\D�0�X�M���r��M��`�h+zY�"v_ �6��¹璀{ڸ̯���w��>YU��m��R���9���*��fnq_
���d���k�+9@;:X�5�����g oV��,�[%��Ϲ�!�dK)GY��N/M
z���h�������?t�4(�h�`\�qC�A���N��=<p8�����O�
����G�P��z�|�I�G��-$�����l������M��Hg�,Aڳ��a;_θ��V�CC��u��G���}�ʵpt �>�>Z�Ɏ@�E�0r̖%�@Q	���L�>��Ë.b��o;��
J���"��)P�"��N.st�}�2�Y��W�1e�J�r+y*~HS%2X�Y���3�5�T�K�f�H�J%8%����RN�X��vA=3���,,D䇈�)�ޭFwsɳ碣�չ��n��J-7�pNWz��W��(8J���ۘ<�x�)�!&DC�f�J��̢L�%'fW)���D�k�I�r�u�#�n�akC�=1�C���r��#�T�r�I�ᮒ�������iEG{n��l.G�DA&�Cp��S�;�X#Ж�7��L�9oJ��k����8Z��f�t�r%�%����3]e
YI��ԛ�h�:?�/u��o�}ѮMv"Te3n�8����P�v��GV=Y�F�d�N[�0_OөU֣���"6�t�AvN;������B������6gX��+��;	+vڴ�XlxVHYEB    6184     f80��w������ �8Z�^9�]��,��M�qQ�C�v�U��ǚTO7����{IhG�]9��\�H��w��p=��h̰�Iw�ݴ����#�a��	��O��DJ����XG^�4RD�O�l�����qFu2B�y�ʑ9�6¾��{e���b9 ��n	���п���5~�9*����c6��&˿
��U�Cۄ8٭a���YV�N�8
����`��~$�876����pw�;�-�����͟�[Y�F8����s7B]�2e�Jg�+W(��!�ψU����PA�k�m���J���3<_�1J�����D���Q�L�MMD¹&���r6�C+*�>�r3�Nme"v��|�ܤ �)�h�{�7ܨt�歠�^PG��>2L�_��W�\���aj��~Z�=�)q�@F���xm���k����E+d
�Z�H%�	��5M<)�����i���5���բVu� u�P���+�3�f���������sF��7�-	�؊��C>ǲΦ4��Juy�T�����WpN�4f���;3�	��R(v�k���T½��'B��n��Or
�;����3�jZ���n!xd��'�.�=�ǔ�cQ����_PMN��}pܞL��gqJ$�/+[�����(�7ʲ�E��BmG�0ʾ��[�e[����
�i(�Z� �+n�ÖtU>iL7��υZ����5��
]�ӂ��"Z$�~A,@�9���2����gu���C���اg���i��ҔpV����I�o~�]�}�̑YK�,���2��������sL��V{��!��f�����8��+���,������"��M����,�M~{&1��0o�����L�'�/%��g�cLP��S�d��ri��O�ξ�cj\�Z5�j/�R��Z*Q�t|�}���vW
^�Y��[�ۡ�/>��f{짰�Z?��f����@�TCI�"XC��s/O
���#s)������E=A���*�Љ�u*�437�'��tAn�ٽ�U����?<��_^���w���oZ��AS"���`�|��g�f�!{:�1�:�W�J�s��WAv�o	@��b/������;r�a��#6,�;MV���xd)���	��>~;i�R�����]�2���bl��:0�;��D_�;�A��	s��w�� �^ژ�9[�`���^�Y���2_�>ʃX����h}tխ|ɜ0�b��U��Z�n�.T�S�.[�y 0�iuʲ�迲�
Ҿ@��?i���	ů�[Ê�d�ICN�?t�30ˌ�5�i�]�,<f�Ȋ@d,������U|���{.�ZԎQ���摙�|�N&u^�q����YsM���eR�f�E:$�mZ�����͊HA�d�M���ly����h�kSJ���SI�jb/�L����S^%��ksʢ.�Z��׹j/��O����?k���k}�I�$q0�(s��<������m3��	p>���R����"����@��H/�ֆ��@�+�)Z!{0��[i��#L�}O��0ے
��	�{쌗�r�E4l�>�?��1�o�{��NQ����y�
�{2t�ȕC-�3�Quq��(�'J^Ga��������@���&�g���轥�kMJg~���2z�W�/f�%��c��&��8D����aۡ�,�����B��%�%wU^5�Ȇ������<�	�6��Y��=l�@I���
���>s<����cf%��L����	 �i+��S����F�y��;��Ed1�EHq�o�K+-���C��Z��x��Y���J<�����Ϣ-kc���t�*�3J��k�|,�q�RTȱ����]��-M���l��e*����{��㾀�݁�1p�sx�����4�8klf�q_�z�Lm���h�˺�C�}����+�nĽZ���"����G^�4G��5��k0�G�W1M\���
�	#Tl�F�NSg��Z� b���M���{��~�� |iB)���j�5���z��S���ҟ�����MdQ�[�3A��
T6���#���e���*�%L�/˭�^K�"�PbY��}!�������}�諌R �����%FD8��g���񂺛o��6K{R��ܣ"DHG�w�yP7Axd<T�`8+^H��x���Jm���qE|Z��xI"\�7���a�ռ牰�-tL�@MJ���@#y�����(�&H�Q��_Sv�E�O��]�!+z��Z���w7g��an.�W�&{��w�O#m�3@')��B�W��K�<j�r����!�e#�`b~���Vcn5ۥ1(�k➇L�f=�o5�#!�wEK�ԉ�0����My8jҷړ:շ���ü�4���Aw��g���&Ԭ��/�Xf��
�
,��d����j�N����`v���*�1e^�c�n�%%v��Mv4�R���Hh�&u��{&�A�O�[;b,:�E#pC-c �/�pht�˸�eg�f���h���(e��d���$��{[J�@j�9�驞��f���{��UzQ1Op!8�G�;��S�5��`r4Np�Oy��|
�NJ���#��1�=�n1Rs

OI�3���M}�#���G��t~�-����ā���N4�`<����=���K$l�����ш1⤚ѿ��je��.)�2��X�tc�2�(ҩ^~�s��1ΡH�9��8Z/�:)s��&��ոp���\��K�qU3wC�w<c�T)�8��מ1m	����� �y�/Ty`Q1�H��F�Kt����x(���G��ԫHIL8A��/a���Q���(O�'M4�ɚ�#{�U�c�~�r��tv�_���:�ꬰ]l�����R7�$$��S�&�lj��<���1׎�e�f��V�8�J/��X�@�0`M��{�!u���)8�r��	�M�q�܂L�3}Σ��k�䈈	����w�:��K!6w'	�������`�Yn��H�q��;���z��l�`��Z$���6\��h��#R���aW�ϿJ���>B����[�&��J��� ��`����FC�-��{/��.�t<J��	;��]�
" �#�|�����n`����g�j�?���;���4����;��XϗE�z��H�}㔿��7|W�vp�g�b�Hd�9z8�\pU��{����s�k��j"���a����4����{��\�6��G��=��t膠m��Ot�r^�Dq�v�$��MK��S��:�6V�J���3������:2A����"�`��JTm#tyz�_�+��=���2zn(��Z�_�������k�y��T&� ��"� �v���ɗ��|��k��(K.�ڧ��Q�ݍ�7��ձ{�g�3iA�����uo����V�a�����w�zbV��\�D��G���lh�D:�T���x����j�a�6��k0�/���v>� ��En*�ϭ���}!�����!�<㌳����V (7����=�p~i��~�T2lP$-
<��#\�:YR��^ur|,Ƶ^;3��a	0�'�Irxυ,w�F�SL�f��Ǎ^����Y�S��|�%��6�8���t{�����]���{I4w��� _x�E'۪��?�ifbT��d�X�sC�O[�,���� ����/(	�?�-���3�2�����mK[���~s�&��'�07�o.p��
���);k|���S��=�-I�'ކ�8�ʹ , �jǊ4e��(EI4k�h�AN�֘3�ný��ż�g=>h>�3�:���U6�����89�T!���� �Œj��铫��}R��=~)���f)sj�?�4������/��O���q�m�
)�������.�D:��5�Ɩ�|	i�����