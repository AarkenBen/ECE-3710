XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3�B�����8�c�$xۓ��T����{�C��j��j�V8�(\f��*����u��$�(�g��z�՜ټ�����댖�8�A�&>m�Q�~�s��c����E�` �Q���k7$gT��������E+��jq�d/c����픧��JWT��o9�F@\�׵��>$���GH����ä~�M9=�ڼ�65�~uM�*�����H��G�*���y���D�,��s��Üv}���Q#�;Թ��}�k�,1��O���t�D���l[/����q�P8Y($�*=Qس����}�]b�'�/i���ѣpZ�>`�� m�����y��!Q����YzNKv3����$8$���&����(�"�)�t��d���]��f�����j��*����4EE�Y�{8>�=O�C�6���
�@���J
י���u�.��xl�_G��u̢�7�����>C�w��DFh^)}
}�2��XϊK��S*�����:��;�~�����I�r��Y9	�[����:h�i��Lݱu������8��I*��h��� `Q�||��M,�u�A�]�#p�4��t���jlf�E�ĵK(�c(�b��\b6��G@E�_cԂ��W�6L�w��e��6��I�|p@ ����
,��t���Y���A��۝g@+����Ӈ�a�4~_�=yޭQ�u�Z�p������S�"n��OLI�m�x�z��dN`#���6��\s`�y���>7#��S-�`Q���۽��z��ƚXlxVHYEB    1427     840A��U�o��ֺ���G���XId-�yQ;=>�(OIH� ���p�d�G�>s+՛r�:z2����_����˺,��P�Ȗ�N&7&Eldշ���z����a�����/���5#��� V���7�%�=k���@9Fd��	0$Ԙ����*��n�򊳋6��e�o>��|�{d��M�L�*?�]?��!,8P��gV�,<��#V&��EB!@%7[��5��Knefu!���B���)��'�@YU\KIF�Q���I
�D�����މȷ�;� mg��U�Ɯ�S���[0�7�D��󩥟軭�=Z7�Q�A�]ܴ��"�̰�cg���+�Af?�Ɲ.��yG�M��r�?&�	�Ɗ[� ��}F2L�/�<����aA����Y��Ż�̦�E�̸H���T�t��VP�
�F�ÉӋ�<y�\��qt�^�X��&Eϒ?�j�t�%�U� Zx����liB���	N��M��y����P�� �m�M�f�P���e���[Q���ڇv'y3�yIN��NpUȎ�rު���|{��3�Ԗ
~ڑ�8�M#w(M.���Sf�����xq������#��9�7u~��#�,�JΌ�V�u�$��19!�N�c����p3�iw�7g�ubV�8
�Rlr@YGC�]pP��~&�"��1�t�1!}*^k�%�E��� zv+��L��~<m��2<����.�}�u҄�x��������[���t�}?��n]:M��P.I�@���=������ldme�t�AGfd��,羃O�+G4�UN��}���kD��)�K1A��ͺ���N�����E�}s���`��T�� �6���Pz��Զǚ��t�޺��g���L�)|�6���/8(a�_Nc]���)������p�u�[��>Zc�����_��Ӛw�Z[G�o_灆���ۭpN�o[��w�m���	eܕx��O^)��yMjqcՋ�X�Yl��R���r�(���G�lp��Q�Ss��m���>y�:Z ��-��s�Z�81�~�����*^ro �i�c��bk�ΤE�6h�ȉ@az�Ϭ�AR�4V!m�H��O�5����ت���kF�@
��np��R¶\�!��/3~O>x���%�9�?V���#����Wu�9rU>S��5X�o��}Y��2����H']
�k����a`���Uq��N��Y&Q���xm�Pw���#��P�AQ���j�h$��/5=-y�oUS4%g��m㭭$pB��D)�Gz�](�K�r��[���sg���;�}˯Z����uڎ�j����WO�;���D���U�*�"���X��mG��ּW�-����z�����3Ș�^^�@GCr- ���1��/S-{�����b����p����W�F����F�}Ĩ��#�-z ��h�HԷg	�,��&{�X���Fd�n�S{ݵ���Bd�a�_�g3������ngj^�66��(�8�������)1��x��}gB��2r�`P�/	'�r��H<��^c2XhlE�D��������<e�>���Y�F
��~�V��&��"��l��V���T�����Uo#�[���>x�S�)�Z��"��%���g�D�^���l��Xё��B�\<���lp�!�Ⱦ耧���߭"���=C��r�ѣ��ߏ�w�}�.���#��	�{�ck K��ɿ��^&�9����М�OLn%�7>e�1�����s�%e~`�.��|	��`|���7>����5k�0�=�hz46_����ɛ��:G��u���ƴ�;c�!δ���5��rg.���$)gA��H �^w�P~�+�aw����@�y2�ٽ{݄��Kt��:�4.9Q#|��B-���F[-�,��d����K��cʧ�8%�0��N�K������X4���0L���`1���pK�!�%�x�L��Q|��K]�C:���¨E����se�#y�TLe*C5d#l�/uƫr,%e᭫�����y5T���w��^3����n������U&�����f�^��q)�
U=Lve��8!��)6��Z��