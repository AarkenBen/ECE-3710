XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��jt���[{�cģJ����(5yM����X?;L��E��&��9Ӥ��n���k���Tff��z����wM��#t�,�BC����0�[���(c,�"l�k��|�N�V���k��i㹋2�6B'E�%�H��dO��_�b�Dj`�Ŏ�9=i�_�a�űa�l��r��<�y[x����eX��A�r��r4j��� h�
ڄ'	�[���W�w��:���d�cN��?�F���bTa�b�f��������k��#.E�>����foi��	X�o)
�9ı���vm y�\ؼ���MD$��!>���~ �5=?|ӥ���u�D2O}b�VbV�"`>xח�r����)E��Acz��]_)�cS������|!������,�0�C1�9T��^�������t\ה��~�Yd���roK�$x��O��1:P;	��y_B��L�V�a.�Yj�2��@q���L�{���M[@HĴ}H�M�*��B�������\�[�@wi��c��C�G8�*ח�rݶ����l�����42��L(N-}�tH��3m�_Je�K��uj�Q�:Dg���]-l�Gջ�؇�e*�lU�pC������LX�S����>��h��3�[g"Q�%�'5�(#��Bᗆ�Q��c>�ll���vbKp�F���A��Ә�X �4�!D���ĥG~5N6Qw&�Nw���YB��B]7���Z[H�J���-)� �E2S��=XlxVHYEB    9de1    16703���<�2���ħ�5���e�'��knfm����汫� ��,Q2��r�B���-�L��Й��df�����7�+2�"H%�Q��"bh���}��l�?+��C֔@A�Պy�tg�F8�gs�?���ew	�?�qђVy��A���f�d��mF�S���?���;�E�������H��L`O���7��;`�9 *�������P�vz�o�T,�q-���110E�Q�4��X���=�0���X�V��<Lh��f�0�Y��XW�\|�4�쭺����f�}��?�WM�����s	-�%k���$��q�|�
z�� 9m�ġM['V�֪������.���B�]����ux�<hq�e�~W�t[����trM�:�i?�p���֮m`/���C��5�+�c%{a�^�xז�j\����o�>슗E��)*~ڔ��~�r��3�3���P��Lv,�+ 53ln�����;c�.͟l�?���x�ẋ(?���I7c�6�c�Fؾ�s#'YB�W-�hyZ+��W��qe�+�7�|\�j� �)��d�Ŝ�
7N�����ͫ���,�ʻ��!ގ�`��
||�0%�ʼGJ���M�;A����X�74f���"�+���ԌB+N�@%��c���n���T\D�A��;���}��T*kQ�5!w��.��	��JM��1l�Lw��h8��,J���Ē������΋)[���� vr��(W=:/vT,]5�v�\I
��d��]��B7m-�k�<� �r/����+P��L�eʇ�#%`j���u<TQ>]u���In��֝�d<M�%3�T42��b&ڌL�\�B�NqW�{h�=�a�L�`�M���j7�eJ��zu��t�:lו�d�N][�y�{�@��k����n>�d�MIv�,��4��mۭE�Y-������pϖ{p�Y�����<���켡 �.8��2������!����b���=#̍#��k�N��V�.�/g�$:I�[D�p{_ӻi��#Ό��W#`�j�I�B��C!f��f���z��]pLJ �$Z=�~s&�v�J��C��P�6��=�;��[��d��J/��ﾭ���/P�⏦�X�kϯSQĎ��F!����Ah�9�/�X%5�s*r�,&���"R��)�|��Gl�℩T2��D���i�QM�"�]e���߻���R׹J4?��Ex�3��-�?J<�4�f�U���a�3��ѵY���<�5��l�"��$*f�'?�����CjKc��n@����ͧ�����ߥd��g����i$�
���g���y ���!l���������ʙ��q�$�E��ذ�]���=�,��u�����	�V~vpf�\����3��W���~�9��	T�	X�9�|"�P_���L1)O��N���cV�V�?;�Z�=-S��"�o��b���;��Dg�޾���F�`�_���8<m{<Im)��Q��Ǳ>����Zmk�ҤL��q������P�V~�*!O`��گ�Ը��þ���{�
)v<��n��i@}]N"X�'�>��)Kl�k�LG8��Cm)�h{n�N��v߻!��pw\y鮂�e�xeo�\]KBŊ(���;�ل܁���8��@�K�ã�̂�~|�9D��~,c���%.���1z��<�+�����cS��6�)���j|��Y;hP��j��)�W����_��z��0[�V®�M�����`-Zd[�
"�&/�t��� ��}\n_���0Cn�Q5��vWI{����[|�أ�bu9�,a%�V������1�u�w)<B_�z|�����J��E�$T�̶E&�Peus�Y�;V=l��$%�Q%�ً�Wm�앏p��-S׉��EuyRGU�ͫ{g�1��#�/��3^��]G)������U�Q�>���6���б*��&a�۹muY�}�H:|UW�N�-2���U_}��;�k W�O��a;�>��s=H'�s�BN�Yf����tc�[ �p�n��G3V���΁��o�T�.��>|ѱ��m�����	U�0D6X�[��H1?{��<�γ_�z�� �X�Ԅ$��t+9����k��W�+ud��"nNޝn�> �>��sq!�L��d?��I��57�{>o8�y�N�m�C	��! �ȣGMŊ��f��C&��NE��=V۪\^���� � ��}��̔'\��:�~5�FIڍP���c�d�1�1���k��G�s~�T���;KH��ٙd���L�/���Ǔrk� �!̰���:�/a�� ���"�I4�iD,������X)�����M�V��2��(�C^2��+R�YN8�D>0�p/Ɂ��a�F�ɏ���:[+��C*���~OJ�E�w��4��Ȉ�r4��ԽC���ךkΧ��G�Ӹ2,ȫ�#Q��K��ɪ�,��\P@a�VE�B�8�������T��,$�e��k)=�2��n:�D�C�_f�\q��PO�������]^޼c�����Y�z���dҥV�&tQBMN��p�؜�w:��_'�]_��>�i���? ��A���:��8$�C�����u]i(��3�:�|z��	��ڜ[�nfCg<���,3U���`6�N!*-Hg.Vs������3�mg��s���b��A��fr�,�q9�h~�A��d^$_l�m��	��V�`��o#��yhN&J�"��#.HR�W���y{ ���#ܕ*�߰���<*ݷ�Ee>���0{;��p��f�WV��e���s�ɻ��hv�	nSj�R��I�����-tݯ�L#xm[Jhl��� );n���r��ai��۰�>�Z4��	n�qZ*�>�m;��V	4���.@���F}!�G����[����5�M���c���)C]��Y1�]�6z�O���?��K����pA���t����
�Y�!�e+�����ԍ����W�Mp�Un��j�9����<7��(
���V?Gӟ�7=������1\�MGg�#�դ�G��i�"fOvģ\qp[��ta@�O�/P���aـ����M3g�>��U[��5�z	����7�`����NH6���@��J��3�cx��Z��� ��^^�@��T|��E�u�����
�mU9j�k�m.+�ʙ蝒����@@=�~g7����_�i��޶ׂ
蕽��
U��-"��&&ͻ}��t+���i��'g�O�K���R���S�`J$��'ΫO�Pw0[��V��/��(��4�S� a[�ȥ;� ��Fu!����~l�~�*S(Yv&Z�TP�������F�fB8�kOv�Bj�$��fi��D:m/9
��	�vgO�F>��5=�d�2����`�.����8��tr��N��R~�E݋E����(�F�2�J�!�"�S&�����!��[��*[R9{>�%�V��pg����m'Y�T�p�ݱ�Ϻ\�x<�#5l��l��.FuI+SV����@ G*�\��y[��@|1������ɭ�z��)Jq�?��Ԁ�~�D�(C^MNmf����wbTl��'��06	��M�!��%b�Ӕ��n�pT5�qfnr��~h�RA�<��������X��ҍ�1��0r��D�m.�]��h3*6b"�[�Ϊ�����_���h��q� 1�W'��}O}��筪k��ܠ9Bi���h�U�}��q�έ=Y��Z�qν��~�``���!^��%+"�l�q��`���pwm��� ��l��X5Ғ�|+��,Hʊa鸧>�"���nZa�H����9�"J\n����8o�s�Ԙ���z�-�R���xNU���Hsv����Y�i���,��tޝ��,Ǣ�)�[]�W
F��
E�� ��W{iᙘ��Tm���S)�q�e-n.V(#7�UB���.�� +��Vxt�f�FARtT�ځ���^�)�.��;ro�2�	���SAdf���J>6���UOkhG>�z�g�������oƥn�+�$�,�Ҿ��,�Y��ی�,���^�!�\���*��6���Vg�)@����4W�!���Q��B=}�KY)[����fJۀ6��	[��������<����i�q���/�N��bv�x(z���!�r�G]_�/y��0��_sW�^�a��u��yE��q׉!�ОY!�G/y��l��n�f�t_~&��y����a�y��T�N �������42�h�Фp�L����(>�V�E��O��w�)���l���G�]����L�}Yi��>��\/�_�r���&���V�}cj�UkcA�;���o�]Tz섻�X�x��ݚ>ْ�������J˛���
��<��Coڤc�����������4w��6LeZ�I1a�F�6��B1�H��>��ٙ�)@(9�3k���S���Ðh������M���Q�a�����76o�.c$z�2&>�N7w��y�G�|8�?Ɓ��J�;�<o��5�ō�;�\������@i��#Ag����o�H�
Xv�(�:�Ė���[)����ۛ�QR,b'�o݄���ǧ��&���2��Z���R~��_ cZ�h.,�-Tc�=B���ɹ�Z'ܡ&�9�g0�L�%�F���&��\&��������x�ŵh��{�����N��	X0�6T��Y,c[@��Fc�� 3��?9񳏠�~0�sC���}E����ƌ��5 o�<:�NS}_�e��9��"f�"8� C�i�i��p���>�+-NC��*��M,x'����p�"&=VL>�� �F\P�0��¨��r�b�՞��8�X�p����#
r��%�!]��<�:���3�����ܯ���v������0߱%J�������h�,'=��3v���W��	X�lcī��M�����;Yq�I����߰�Y�8�)�B8粮0`>���m���v�O5�*%�-q�MD;pzG�"����e���m��� �i]h���Hh�7�-ȿ�L=���[�gbn[.t<A�T��7ʌ�������#�W+�]����O�2i29f�����Y9�R8���}�EI�m�>����eGS��I��A���&�󪵃D5OnNV���&��e-��zwߋ��7jS*���\��R�z�2���O����x/�|J]�d�3:�uϥE��m����:��[�Jڭ��Ϛ�-��e7��`3r���6�LBEfZ@m����9]T�@����?X�m�����˼��J�oI��5*㗒jo��#���jDg��D5�eKë�ɿ�B�dH �e���V˳w��Chm���&�9�3ϰ)3[?�h�>���ƕ�$�!]�~�k�翕9`�����k��/#:,�-�ԛ�e�7�\H�Ql>s��՞�?��HC�$X�&�b�D��m��(�|T��ÒA���G[
�w�a
�����a�n=@vq|w��kw]vU,�%���_��n�'�ujM����e�����5��o���&B�lݓ`��{U��/�$��aB�q��wO_�3}�xm����OR����֟����p�Q�8�{��AZ�����os]�Pܦ�5�