XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�3��2>��x��|���r�=�B�N����,���˝��V�vo��,���I����ߑ��`/w~�T5R�|��C��-p�Z�3�*�#1��C���b��v���	g���G���A�ք(��X��v�u���8H oK�� �+�!���=���wҰՙ]�7�s���|�X�=	J7ׅ�d��\��"���a������h�N���B:����\/t/
%�߶X{�&�}i���G���������܂( I��A~�}��� �����C��k�k<�����V�{?)�p'l4�,��-��u�zy栦�8�	�F�������z�2[3� ��+=EhC4�\yס����:$��b�s@�&�/���D�\���z��e�Mvr���z^_@R�*+q�c'QѨ��*^MFAM����W(v��w��WpW���ä-Qtx��*ϑ�Z���P=�3��J�40��ou1)�M����-n��C4�\�O~L���A��'��@؊��Jߡ�xD�S�O�����"�[�9�M���t����0��������l;�j(�Rj;�c�K���H1�h�Z2H����xp������_���Y�8��4���7��*����W������k {�1���u����6���R��J�.���?l��&�_M:���,Wn;	�w��OY��w<gv�`�ΰA�N���d�f�ݏ���X���̦ u&_�1bJ<-��bJ�'uxw�XlxVHYEB    9732    14d0�ko���X������:�\#T �?O��+��)K����<����5����V������<�@X��!e�Xs��0痚F��u�3d;t��)`(4h� �k�W��T#��!D�� �HN]Սi���W�KT�縒�P���/���M���ݑ=� r�P�61X1|)����.y��RLlz��<A�o7��:�(�u ��ܩc��������ơ�ƍ�����&�+�����*�dk�]^���X�2�%�͔�$��}��H�o-�_��O(��f���à���2��N��6M���P��q�lj�a��@�N�嫍p���j�TI7�x�U5��?A;��S��<�7�D�8���ȋ��<s�N~�D����h�h���zm,h��wD$��C�Ӱ1nq�:,���(�G���$I�H'I�����%Y%G�w�##A��^j��^�a�u�����V,�����h�`��+�t�w��JúE����(f ���	���	������,��3vn�X���`���=��`�3�5,5���b�Pˣ�}&��lz�Ϝi��(�M$3����,D�%��7"�I,�GT��u������o���5�cs��c���/�t]�6s��XNd	�Q�T�E��L��S���.$�9�� �U%����(�^����Z�O���ci^�Y~G�(<tOu�ߠ8��c��hW��N�/�)}��M��ܝbS�'38 ���8l��[%�w�~�v?=���"m�G�س@�_�0=b�������6�5�l�~d��Ab7s+����2����J�.A�2��TqR�ƫ���������;�j���6��E��������I�k��#7Y��W'�n�RXC���z�}6_��ރ9 �V��>[ �A*��J�㖣�B2���.IE������}I����p��	gr��.�E��ɣ�-�s��Hu?��K^����XH�%v�̕jh����,W)���I�݅�>�-�ŗ|�\��������������C.��st��48ӡ��׭���H&�#��~����S����t&�o� ,��ֻ��Q��ӌ�5 [S��%��څm�d|�*����d4S��{��.Ή|��K]�NH��^�Q�&\M�c�	�ѓN/j�:8.:���-�<lݖ�9۔��ށ��9WW=���3T�4������D���N��#H��;�/�wW6u��`LM�T�@\٬�����Xxi���S �xH`<����D�ƪ��<B�\�k�3��K��F|�[}���i�n�g2P֤$VK�`o��Vw��ˌʜ�˽�X�� F�?��T�[̭��L� rC�,4Zká"������؄c����OB��k�w�WP��;l�B��?c��J�x�P4��*R}i��������?@.#�C6*����=��1��׀DX��y�@1Ս���|%�;MZ2�։2Ļ�@�A��\i~�|�k)��nG�
(�7:�j
{V{�_�����ӏ����C��p�����Z��ld��h�����FoG��3��JOP�ϖ�s�ܖ����5�q66?ضFU�;�3ϯn׹�Ʒ���`���i>���ԑ3lt�ӹ����0�cً��6r5��~�/��@�9ˁ�����@65�|�B&��|��Y�i�(h���8$R�REUĄE߀ߑX��I��*��G��F�._�,�T�7�.
�X�O�$�Em:�=#�p�˽� ��o{�-���׏?� `	�tHuM����p\H��u
ʈ4>`��>�ͩ� ݨ���<���!��[F��P��B�-!�E[���-��V	��Pߤ��$3*���̂�߯�U"���m�1�VJZz���S��4+��5��"+/6S�R(�����D
���^ɫ�@lL�KA��-���@��w�� �� �՜/��|���=��d<Y�,��PY{������}"��
�r����d���Ν�P�N��x�G���"w���}:^*�����/a�YT�Y�!�A﹡������	�����7.�uu�>��HԼ1��>���y�,�����4e�m�ĥc�d��$�:�G����}��W�ԇ+}K��F:ݣ^�x~�!�]�3�����|e8]��]oz�E3:���K������,���󠢴�ߤ+�[�04�C����3^+��l�&_��q������a)(~��uÛv�5ɾz����˱��M�s�Bi�@E��z��j~o��������a�x ���1�X�ǒJg��e���s8�@Hr�h�&����DZ#Kq��Y�7�BA���1�a��B�u(���P&�<�&;{�iV�P�0���z����%�v�c���U[A��@ՙ�ƙ@N���Z�9����wLSu��!1���v�vF�y4��8���X��+ȂC{�d������<|j�
��G��GD�s,�I"��sfO�tT�@"��&�o��X�����8s���m1����'�#���؍���w��=KP�n}�f�wy�oB�����P��mme��D�Rá���n�y����!"���A��|vY2�Y凌��B1�ˑ�.�mF�G7�����O�4ʥ�j�H,�ߋR��K�w߄�o�C�ji�7' B 2�*�=�cW��P����|�ە��L>1d�����jް[��yX���_B�V���)v�ą;�T5y	7���C= �O������' �B�;r&R�M��g�
߄:�]UJSh.>.t �<��8�i��vp��Q(��TK��9k�_��)�1���dY%�Z쉉����kh!N�౛��K,��{�i�ޣ�Kޤ�&
޻�Q�A��1��H�Q��{�;�&J襻���a�ٷ��$�ם���a&�'�rj���4��$�±�3 I{���q���:`�U̝"p>g �M�3�� ��L�_842b��@����N��_@J�yk϶aЄ7���J� ���cҞ��O%��Byf6��LAbقIA�y99X�2i���]�F�5sI,��*�y�/8ˀ&����Z�.j��n�����Z_��Ӯ�Rp�|�,��y�5��[k5#�敌r��BF�M�����������_ϱ�
,����1� ���G��N���L���
B{2��@�k/OS@-7�`�>�>��z��.YCS�R�,x�7��*���_�~%jo�v��p�B��ߓ�s�!o�"Ї$[����+�m�� =������,�x��,9�W�r�#�9��6�ј]�����~}M�4 ����X`�S~g��4���>}��Î�$�L�����ߙ#+�t�D���z'`v�5����V��VQ���@gΰN6PBKD�;&\�zˤT��d��F��4�v�q^��G	�rpŐ�U�@%�I����`eҗ�QrJ�2��V���D�}ՖnQ�Z���Qϥ+�KȒ�ZLW���(��}C��$�8��ͳP����tW<"�;���ru	!�#YD��:<�^(��E���Lt���{�qC ��#���&};��.y����n�lY�_��N��+�
Y]W���p����S�B��C���Fm6LJ���Ċ��X�Ķ����G���gg�0Έ��Z�[�0��5�Yv�x�PΛ�5d��SNỲ9Py�!W��l�I���{tx[�5�A*`�tA�>�xH�V��K��k��JY#vD�g�Esoo6��?c  [}Ð�`��IPjt�Ǆ�v@�O[�Or��� ?����L��
I��{��eț�m�-��/��M�`'�#����i	�%��
R
�]A�2��5��oW�������d���ň� ��Y!帳Դ������x{Zv��^ӧMs��dQ9��X	�J36F�\-��W��}��7ϼi�ǹ\�{�i9�ŕn=@�&���B�����MX5]י�W�rN��巇�7`9���|��e��!��ӧr17�-6G�-�H+I�z_��0,�z� Q�D��h�>5���(�ل�x�`{�aOПme�y�K��<��� F3!�l���We��>�J�a�O +U&��_J<��i�C\�Q.AAh�@�;�Wi�����8)��5^�y�W�Yƞ�v�}�	�H�u+Qor�G�J�����Z��0]� ����!��<v���� �������M,�C/�,���Wq���.1��������)�k�ѧ���H�r� ��t]����������rA�d�@��o1t��:����*�{jUR�U}��OׯG岾����V�XZ��]HK�5�]
�=��0�M6���E����$'��cBV���+����
9{��}�z�Is.���I�?���̜�������ؐ�"����𫫜u\7vrЖ̘��7L22���(��2�(�o �W��EJw ��v6����ј����l��/�/!xN+�H��B���4G��:���拮�VE�� �Q�h�!��:���r�Zdu�5;��gy��=yL�z��&����ҧ���;�����f<7mw����og �+�ܱЊ�?��^Q?����t_�mZK�=
㫏)36H¢��1.�'��tH�~�Q/)�����#�[���vf<$$�4��&���O�(���W���/��^�e�
���x��\��X�˜���u�\��U{�:[S-�5�Ɵ��7���b�H�Mh`k2 3a
]i�ƛQ��ᖍ�y�a��U�
v0/�3<���B��@i�k�뺙��U�~FKi���V"�x'�Ol��vm���;ӄO]�����Ѳ��Ta���K��-��ڿbS�N��W��h�:&z���}�N������Ըr�$�⫹�۪߼��~*&���B��KFu��JZ��3Y��^:/��]��:hh�5�g�4[`ZFŔ��:}Ax<'d�)JX¶�}�����rX�Ϙ�O����")K)�z;��s/��V��2^�����wA�޻���7.2\�Q�lp�k�n@A�!}ws;G_.���®�	r΍�Խh���<�٧@n��8Ȁ8��'���jjس�H�#��>��JD�]�V��\��Ι&��d�˪�Sc_��C���(<���p�`L����*�e����:�!���v�������2��F%;�V}J�kҳ�X�k���!~� �ŷ胊�=c�^W)��ނw��$vs�&���� �6�����h�Vߕ�G�5g�����=��T�ÎVw)}���s�&���~���