XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q~���K�+���|�g�n�������YBqH�A���aJהa�6�^�� �}|U������A�zwL��l>�_��k,��мO�r++�F}��n���@1C�%L�Tq;2�m4�\��5��"��g���eK�n2\�as�Tp*�5��P�@b5��g��|��!C��Y�pТ�<9���s����~N伙� ��o�p��+�
�m�Ba
��TpՍC;LGf��6t;t�z�<��@p9k4�{�ʵny@g��5p�~݅Y���rH�[�Fx����4�g�ro�����P�:z��W~�W��i��b�^x�
��&���n'W�HI��D;�:ǫm*YD��7�Kz���I�ؕ�>��=���^rɘ��X��ɦ�?81�
���ө}'��w�QcR��)Ԇ��HB��ؑ|^������r�+�P�� �Z�d�2���Cᐾ�3������ ��5gl���R�LD���Ȳ�>��N|����G4�IFw9�,Dڶ t���|���Pt�8�I{��w�Jm�xL�y�b.���D�2�q˨�*�$����� ����c�f�/��
c�D�gTS���Wu}�{5����H"oV¤`L��h0�YT�U�H�IB�k�c"�*���H�[7��l";�⽓	�4�֛D S�ˣ��<
%�QFa�#�1\�����.f�(``UK��{��+-����U��t}�I�%~~�A:�N'�&4���@��ժR��'sY\U���K8���0�XlxVHYEB    2e55     b00�� #��L�J=��r��s�^@'��k�q9���:1|b�����)L�.�m#�ǁ2�j��ٷ��<N�q7@�Zl4'ϩ�/��H���׺�����R���"�KU}���p�����{��W�����f���F&K���m̹� �}j���v ͍}����CkqO���w[C0���l�z��h@�l-��Ǆ��`�`��&���is��bǧ�U����^t}�$><Ц�ܮ,��[����֖iu�xd��ܔ�+5}Y9�'ik�M@;�4����YS�ٓ�$,���"=�Q��v{Q%覮)6��0�Tb�J"��F#ާ.�$0��Y�E�����^����++i����#p��0�p��Ҥ��Tw.�2&�������Q�V�O<���,�9�:�3�ڹ;΁�U��;1=y̒������Xd���~���kү��{ ��3�,��]k��U��^��(��5J��+[�^iW��Z9��5�M����7��g:�2��m޵�ꘃ6���v��V7�D�]%�,q�x������l1��U�l����(آ�f�0����^>�/ҍZ��8I]�.-�/�a}��
��C���v6�k���W~�^�n�������hջ� ����pɎU�Rk=Y;{:�$v1���V�5����<�G�@O�Z��~x�Ez��#>o��2=��O�{'*m���q��X5�k_��Ǻ�ڐl�	�.NS��j�0z�XM<��(Kf������=��e�-w~ˁ.��>Z������p���Ge"(�rz�T�N�/ps9������t�]�a��^�(��>6?p�
T��y@ۏ��b��a<>���]�FgD�{L�3y�#���y�V���:B	�P�qV^LK��37���<O/q�kvJV�m�OU������]��.i����zس� 6
�$�{�XI`L�1QGG��N���ŒK�*��ђw��C����B��y<���6\�P��:KP��u��Xȃ#!a��$�n�R�0Va�����$_enӵ�}�EX��q(�+F�s���oQ�O�o�5���[ހ6Q��Q���
#!�e���)@�΋7E���륀��@�O��I�fR�n�'���ҿ)C�! di<(~��)��3��"#�9c>!W�%��i��λ��_�̆p/�U��x��z��XN��]@�Ȇ�\ �!բI5�J-��0<�&�mz�u�rG���-��6��k�*L�hI�M�T"A^U�`����I�y�.�g����h!�W��󮏮���:J�-51A���@�H��J�e�Nmڄ��sw���bUL�΄��_�'��������9�=�iGfn���b�k6�6�7r�āJ�;iޡ�+��,�aZ��ʐ�hVЬ4h��a�T(��\ۆ�!aL�b���6�F&Eyb���]�N���k$�H"`u�C\i�+�m�6�wZK�'9q�˺aQ�$s�;C��l]Z��_U�@d���s�/GLZߙ9E����j�x*ez�$#�V���:��'Q���cU���Ύ���t�0���5�;����dP8��;��s7�W����s���0ts�ʟ��e�(�~`����z�T+�����.�Tr�Ē�����nΦ�Q6����I�uo�)�j�$���Lc�6���9L������ s�'�	n#��0`������b���"�Y*��s�Wg����|����%+��L�6C��'}��]�%O��d��T*E]���7[�F�# Uf3�f@3�
"�i1��ȩNu�c� �����,��c��9|O)l%�xSa�^�ȇP�7��2l���ƉP!��b�]l]�M0+(&L���;�-�� 1�#��7��@�C�@U���2�8�T��h	�/���8��o�?�#�V���]Kin�ח;fR��v-�b��f��\�X�`���튎V��\E�~\R�CN��Iida�Fz&�\�ܬ�1�n+�n�K�!x�<��[�I��b����86��g"]Ҍj$�Z�o�r����k�J�w>qs�B���$����ȪA�#�p�s�E��k�>}��Y`ݹ�i��Q�_�C�Ij�7Z�_v�PU�\"|� ل�|�(/��H�䊓s4^��$�w��و�lО~G>�j�bPI4ϡ,�@f��¹4�M���=Q'���z�3&�W�L܌�����mn����l�ms�D��e&E��2��l����i���nY��7�]��u���1j�nC~
��z�3��qp�hV�sR�{�Uu��vt���+�І���HS>D�S��	��zՙ*�=wf��KujٵctSβڙ��(���z���WY�%qQ�6�-�e����w~����W�Fư�!�)���9#鶘��?V���!lHPo�>n�K��w�9�� �UE�����Gчo��V��d� �w �p�����P'*\�J6<�f�aLׄ����o=c��f�w�}�`i/u��öA��4[��:S_?<Cq>t�*�/r�_yV���QK̭g�y��f�sh2�o���p�x�0Ų��pT�*ϋ�ת�`��\�ur����H���<Z~!8U=���ZGwU��_1A1����sGL�F��B]�<D�3����ë֮�`�80�(�X3���	�(� ���{@����(��!�D��N���^H寉i޷���'��r�Jm;�|�$��Dn7&�^�T01X��qq/�:�Ly\�� i]����痢h.����?�G�k�s�ɰ�g�&�C�<VV�