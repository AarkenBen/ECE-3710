XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�(te��H�xǍ�T�"�Q���g���-" ��u�pN7L.����u�*c���֕qσ�M����*[�x�a"��n���2�p���4�Yu�^)<v^�Ʈ�H��SB���@Q����p�Ǹ%�w���V7�)�J���۝7�6T�/Ih2��{�����&��x�gC�drc����.�������c4�8q�h��t�֮�3�)��M1B@���B�KR�n��G�M�j�I��f��RZ�K�:�ݛ��5�h~���zh|�0�=��^7��W\;"�歜w֢R�6έ82��rW��g��Y��Hu��.��ǃ�JP��8����׈b�ZV��+Xo���Ld5�N��Â�����/7���nʖ指�B�P,�IES��Ч ^�,T�=C|G�J�3�	���7ϛ�k�V����G�I�o�m�Wr������nsJEa�j���k��m�~�<[	��q��]%ld]ީ<���rJER��-�;Ӽ�Q��3�l ;HC��~-��c��DDP��7~?e��\��űT�:F�wQ�|rW���UZ�������o�>B��Wω\֡j]�
?xx�˻�t�boI��N�*I,��!ž�z�Բ�#�����j�jG'�j���C��Y�X��� J"��٪��YЏ���ic����k$dx���O�vnW
�C�r���vbIL���a�u���z��[�	�������\W�&�D6۰tZY5FeB]�d��݅hjl��
XlxVHYEB    aa52    13d0��px�k�{m�C6v�H��q��YV|�X�6D8���dĞ����������8DN�	�\��Um�I�/�4x&�DO��5��T<8�
��
CӐ�d�*��r��� ��]��y��>��++���*@R��asg>�qT��l'R�)Ka���2�:m��$�1U�]�t�~��]i:^����G��gT�T!��ӞDc�m�
��Զ߭�nq���ҭ��]$�:`�P+��Y0�se�*v�e�����ډ�>R����k�/�8�VŌ�on4|�VC��O%.߮hW����o<���)GML���@Z���`�B���6���-3{����Ǹ�*_T��b�ģ�BN��h�D����.��M������<;�V������D��<of�@��l,��_��*x|;�l̊4|���>�+
�6 ��Ȅ�}D���lxta�0I��籘�B�t���	�����x-
����.�Zq�c��5���''s8�CFVH�utʁ���3���	��(�A�.;s~���yاH��$��@��\;b�M�����Ef�!z�
�W��Ǉ���w��}o��۲:'���~o��.���i�R�$<{�osP�ZOc�Uvo��@ׅR��ةQ$Z*�]h�B���䳗=��#���Ϩ���l�w_fq��rs8\0^V��=�o�Y�?V<[�������4�͛�vcĤ_=�5����י?�_\�Pn�Q��e�@AFm�� FH*��ș�� �����;=ӲuR����x�Zj�\����ΐ��4��: EZ�cb	���6�ܩ�/����Gq9N�cOk��9i�ߕ�ۤXzqv��4a$Mͭ��eyS �6�(��gj��ߚ���Yq�����Ξ���u˞�p�i��Hu�gP�f��I�*���jPa�O��P�o��fuP�f���2���8:�9�_�����T�o��?�;d?��l�`�K��Z��H"�8�F�J������t�!�K"ŰzEp_.�(6�
����n�� &\��,�F(ꐹ���g���W�B�V��%u�U�d�!�O2�h,N;�"�ܘ�@ތ�U��p��n}�j�c<��^f]�9�򥫩�$�*ޟ�i��2�����KҸěٟ&�����G�lrV��pO%�bj�����'1S#m��94#��H�SS�o�"�w��Gĝ�c�c���g�u�P�fK�b�������Gr�Yڎ��m�Soc�!����� ���TO�t����ԯ��-ܒ$���0�Q�T�= kV>)�I�Gz){r�N}cS��i�A�@�e���8����^ SI2I|�D�#	���0��Xn��G��|��8C��� �Ua�b�a�k�	iz_hm��`���/��ɳ k�S��Pz,��Q�Ydz��˺�n���:���6ˤ�^ _ٺ���K��,D�]�Ҩ�l�����)oi�q��|Sֶް��,�W�g?z���''G���P=���\�<��&� �h���B�:�.},� �Xj�{g�f�ǃ5lHZ\�b�X���9T�֢]��5h�A(����g�
Lu�eӨH!_�sa���[��!)�ǡ�� �t'���ϵ��9�ЗyZ�Β��kS�
H�mM��֧���vzB�0�ɵ�Zd�p�Cq&��U*WՅ�h����ap%b��*�?�ĝ��s��J��J�Z��[�b�:�un�ܴ�]ft)��d����Z������m��m&Xa�o�p��5��(_��A|�p�����x��E��)���Mʢ�d����.���t�B�f\��O�� A9�kAd�k8{
��`��懭(�a�����\��=��x���[�-��/
_���o=���CZ�҇ٚt#4��a䞲��"��D9����zaE&ec� x�	�#�3 �BTh��Cm�F��t��7I�]�y�F���]dCS���B�Ň��|�tv`���`H2>�Y��Q��0�z<J���]ݺ�2�C()���N�䑋�)(��S�[��d�11}$�Jŧ쳚�#�	2p�P�E��t`�-�{��u	����Nٍ>��'���cˀ�%�aq��e0^�Ab�ĿT X0�AAH�uͬ��hߕ��5ߤ]{��A_`Y�¹?^͘���L��%
:O�]��������5}h�B�[���*�`p���]q8Bj�b~3��#�m��ѩ��wK��:��CD`�/2����y�Ǎ��������u����q�^y�56�"���0��;p(����矠��ѧo4A�{�c��X2�컳��	Q]��2�y|t�J���*G���q��  BBj�< �NI���Jt��F���]57�e����9<'���"F��7�&�]>���7VD�C��������P�ѽ�@��a���9��ӄ���vf+�3�w仙O5p��������
��@A�4���J��Cˍj�����1}TǕ�/���``K������$.� ���Z����3�h�Us�-��m��ǎ�d��u��q��\���I��Ӯ�bm��W�v}fA�p N>��U��
auJ��˹��ݦ<Ѽ`��h`p��*���f��@PJ3{h5�.A�˥J���AY뵲�YIw��D��K��!8.qJ��":����Z3�r�1��}#��<A����ON1x�ٲ2jV�H*�W�̇� E����	Cޞ�2�OMi}<�AW�Uh�uGkt<���fs��`Ԝ�Hi�Vƥ�J�)PcFnW�D&@�]E���?����D�O��{x,ܙ����*KUo��(#%Tici�j)�d����K}�`1Å?GN-q��2 ��狓��W�)b� �
��S9��Iw3Ƹ`3�ؒ��p�m�U3���8�9��C��L�Q<����������|_O��T������QʒQ�O�F0�5g�D���g�#�����Ɉ�c�	��[�����7���'�!7�����ZT��s��a��b!�l6J�:)���~D��T��>s�%����@kIM��hC<3�H�O�&�T� 83nʚ�Çi�S���^Vcm�g������o�]�|�m�I�2�$a�y-���{`!��[�	�Ew���m�21ȥf ��@=���$I˅���kuP%��'	r����_��
�&i���D�~�5;A��{
�1f�|�	l��>�}��ƴԗE��{�R�"�4�c�6ݛ+�r����.�/">�NJ�$V�����.�L��p�v�S���euL��ŖX�G��W]�*��H�^��1Qw����-q�(ë��y�r� �?�T�a��\��G����Q�����#Bv��P�.H?jc�o�W%��m�nr2���A�>ˏ�q��H�X=��$��-���%��м]%���@�r�X�c��A��$Srd��X+^ G�@i�����2�b�o�r��t�I�S��^�ǂ4haV\�z�-����yqs��?��5�~�Hg�?t�	s�X��Z��V�)�њ��vz��=��f3�v]�͈q�j�*=<�6 V�Ր��n0�FT+��:��Y���W<n�e�c�,� 5��`J��W�a�<8�ȶ���R?�:DW�
�ٔ:_d;��0��g'�|�8���������'�B6!P��=�W������=��E�7 �F�(9�>�ء��HxiD��������Wo�R4��)M���%T��m�$��pPEk�υ!�+���37�:9J�q>X�sWr@W��^�{ђ�}�UE�-�g����9)�e��]� ~9
����X�{�%p���>�dGD�
оu;NdH�������e /TP�R�mM)���X�9!��h����.T��)Φ��z�:����wc��_�
Ȍ�H������^�@8��ԏ�-6B9�̇ȃn���J�G����eq�3�\ܘ��Us�o��$��n�p*�ě��ɼ�:��*Dg�������D��a��4�n!�H����޺8�s y��P��:�R+�|��.�G���[���A�Y�:�����v[�)Wx��;�A.Fo'��E$���ćs{�2d��݅��@.��v�yӨ1b�UZuf���5
 ����.ͻ���؀�eV�,0��!6�C��HZ���HK��_sL�������C&&��󟛾7?l�>�_%�(t�	K���{*��K�3�3f��֯ڜJݝmP���-�!j9��hJ�(�Q1���p�PS�K�$�����q�~�J���lt����2�v�� �iw�I�qhC�W��׏������َ_�8f�(r����(�Ө����0��׋�,Ӏ����C�Ma�D��-���^����G��VY���T�L�-п#Z�椨sCގ��v��s3s@	���I?�s
7����f3�b�� s�2?�Ɣ����.���yC4�6��������E�&���4�ʀ�k�YJ�$JO�j��$
���
�CS�W�"����î��K��qX:���~eqs����z�8v�vE��W[Қ~4�����_ޜ��f�������f�0ԛ�̭-��<ek�^�k��u�8�J-yl��=r�˼q�?��8M�������OR��5�!��!ϥdP��PL,�N����wuL��b�\���ٺW�����M�N�~�.�	xq���]�,�o��~��~W+:���b�,��
��8i�&S�0n�J�[��0����.���w'������[սv[�0Ǧ�BB��<p�Z��;���w|� �%f�E[�ϮfɅf��O�5�Z�!U3�~v�@��!�7�<��ʀ��K�B��Q�����_�,�
��*!�p���=
�X�0��wd��z�����ٗ�ʪP����*پ�$h��Yn�L�}�M���2�k�~!�$�����*����	w���>;FpgQ�
O"��층ҋ<_���Dk��4ܞ`��P�pKn$!��܆�