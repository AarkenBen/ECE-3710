`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:26:59 10/26/2017 
// Design Name: 
// Module Name:    core 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module core(	input clk,

				input[15:0] mem_out,
				input[7:0] servo_in,
				input[7:0] ir_in,
				output[23:0] mem_addr,
				output[7:0] ir_out,
				output[7:0] servo_out,




    		);


endmodule
