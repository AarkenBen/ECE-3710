XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����--s{�*<�Շ>g��ݏ�r��a�&�f��diS���/Y� �mؼ�a��3�Z�����G��s!�FI�Q�P��w�o�"��Y���S�O �hW�j(�h���6�7��`&8b���y�LT���8r��SD#�\ދvwœ�E~z�p�k9�,��b.͞S����xb��y�X���am�l����e���G��\��:v���F�;ErU,DP; o�/����pCF�ɘ�m]���V�o���KֹAgİ ,�����g]�>������q�Y}r}���toILY�]��R�؀�m�u���f���Pw����R�/[�/�hyqP-�=(?�Y�/�}o�57��{%��e����~,��j�r
���`p�k�G���٠[Ӌ��E�՟7�l��bN_&r)L�� ��~ ��I=n
�/1��F}Ws����2}B���A_���	Nn��E����ߦ����Z�Bo�Y��ڻK�f|�c��?O�L�o��n�K�\�D�#$>	TLMBQRE�q7�B5�U6���r���P�DB��ʅ�
����I�,UE��c����c����
À�pM���w�$���ǿ@�����h �H�'շ%7m�����:iߡ��%�y����J<�?��������n�u�����DV����Ց��-޵��)�
A�T��u�k��l��tM�n��~��a;���O�꿄=��ߨ3����9�_��|'���U6����
�D��XlxVHYEB    33bd     c90Gy�1̖��m�G���%���mF��yTLK�����6	y�uq�w�-����OY��&�[;U�{�f\�s���7�E�Y�K�U��P�C��RF��Qz�m������P�z���UZ�쟥)]���#,���6�R�6�k�E�?���)dZ<C�-���d��-�um+��LX{����l���`AxP���XS�p:�6�9������L�a�L~�
9uv�� ��e0o���tKֆG�&@(Č�7����c���1o�Gl�'EYKx-F݅�W|�����.#>7��`\�(5%�O򌼱l����l���VV6�*Ι!<#��o|܊U�fh���m�1���̾�%(��E�
dt����֢��+ĵt&�+�J��!#{��[�� &�_��ŭ~]��/y[%2&�RM��a��=�aa��K��?����|Z���Kq'�ՙ!>9D��Ձ�� �^�.�
3!D^�~�*��3�Q��ac�(��4L�U�뵟$e3�`\�hN&mN��B��@be�P��c����U��Wx.�@�����a�u��uC�#r7Upu�[�\���<֟�wҼ��^~�=�;�1�� 0��`�����.��Z�FۦvnIq��'��Hĭ��hb52��w��|�4	&� ��n3ER֪�GE���Ѕ'�/ǚ?�����o�XS^��k��Yn�J��3�m���c)$�����|OH��"�]Hz�1��)�,F�_��8kupe���P�G�J�:m��c��M�=7YZ���0�l&���V�&�N]ݒ���^F]�9�	%��*�O��\ݓ
NdMO=��k����x�x���cS	�d�rXHbǘv
�V=���ѵF�� �����k�qɽU�9���A��r���,`l�[�@����uE�X�Z#�]�q�1�wBL�Ʋ�k�x������6��-�Ԓ�;�,�=��������_$v[���6����"Gp���^e���2JM����;QX�%�]����Ħ�~t���{�ve��_�b�#�j��=���A�������	�ou����hƼ������McS,�H��&�ؐ%�Z��v�-0�]�6�!`�#�S��55g�h���� R�\Z ��|��lE��L��}x�t�����?ʝ��.\�	(`����@G׀�_��#�N>Y*��oR��b@K� ��A:DG� �ą WM\>'�@�Ml*s��A�N��	�#ڻ�w>�C�dДY������D�Bt�D�\c锦�v��2�!^Rr�FF֒6�l����~�D޽�Na�J�lL�`A��5�3R\]��D�sqWQ��K��>%铑�-�2I���ok5c*��'pb�����Z��#�c4P�R��Vx����[i��~S�x�Bb�e�����A�Y�.���F��Yr8���G�L�� L��҉r�e�Ȣ�^�w��li��������Q(�����u�>�����0� ���	rmr7�@��ն��g[�.����PS���a���J{L�]Q��I�h
6�R�-��_����R
+]X����SQ�;n���!�y��~W������ �	&�.�
�Hݻ�:�ݷ0��i�u������=��'%E�ބ��!CĠ-ç$#����܁r��EN���J~���g&JzA�N�yaǝ�B~��}�f3�pI0	�R�CjE��:�,h(m��q�s�oS�U���?�=6r���94��t�.M'�Lwx,�@<��OlH��YvYU�'u�[�^KE��(��ߺ�d���kg��p�~��Ff��!Q\x��tH�����#���JhE�?W�{�,�����Ƒ���[�u�ĸ�eZ�x�(/Ѳ&�`�u���8�$b	��A0�A�A�F`��r@�V����	?כ��]�x��[H���:5Ȧ3gz�I�t�o'�* �!���u�&�E�2DB;]1�\:�kY��̎L9��TZ.��v�#$8����O�����4�g��F�J&�Z�������	��?�F����[��.�ٹ��BE�~}����F�t��sw������I4��co-��#Y�lK�vbnW4XUQ���*g��^S��m�Δ�h����v���<TQ�-!���!�aw�&4�j��ǻ�kH�܆	J�\����
@����������Շ?�F�X}~_|�Ps,*72��t�z*6My��"P|}����ר>���z9�&��)������O̷�K��ం�5xq]y��(����9�F���>)ܽ�y�C*��YT�OLu3o�Yy�٪89�=��Q�1�A�O,���b��^f^f� =�HC��5�J>��Q�.��D��p �TX�b0O��v��h�p���zi���eñ�>.�^� �*��"�6�Z���h*�G_�7{�Iy ���=�V�Kl@��p���=%�n3���y�Xhuc�:���j��t�:�'̣�Q��b�&I�D3���vb���f<	���J�8~�ñG�s6_Iḃ�*C���^�_�2����[�n�P3�?R�/1 v�|I�&/����*n&s4K�!���\J2�I[tė��m��݀T�bo_�����l|�`��F."�D�tJ���숾�sCsi�:�=�Oώ�8���~F�m�w�+$zQ>��%J0f���������v:HÜv8d*-'�0�fB�ɞ�8w�t�Џy/JKP� E��h� ���e�j��|a�5�>Ѣ["� ��+S�K-��h���<Y��^{��df����|6c+m;4��7� o!��|�E?�+�V�5p;0U�lX� �]Ӑ	Ʉ,!�[��qi��?Y�⪥��ѳ�'�I�6��X��k��=�Q�����؇��w휦� �G gBsÆ&o8;FtԢ���Ξ������(8�PQ�Q�Pl��<`do��N4��ua��#�t.�d,]�=�}+n�!t�NfE����ކk�_�`�tr@�<]z���5��"���q�	��|ό$g1�I��^�G7��:�ԏm��v$(W��h�C��1Uv?����5k#&5��3�rhi�?����W��Q��2o�Qi�e�/�K�f��[�U�Ѽw���-� �x�h!"��'�&��j�e�$V=+g��ڕH�k٪��#gW<tGN�,'