XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[���O&q����v,z@�*�D�#��q,B;�A>�4& [Y&c9�B�`�6�[~��;%Z;�hx�9� ��;��$��Wt}hb����b�A�]��������,�>�o,���|���&+��jX00{Q��&�̦9Q)����0�ci��V��f�}Mp��	��j��k�|V�OP1v	4T��Ũ��.���̻�0��$4=:$�$.q������C���Q2�hLY�Qͣe���/��*����\"0V��)*���R�C�"�(�w'���YGF�lO�#vJث���ަfh1�L>(=RBv��������{�z��|����)���!D!��zG_�A�Ƶ�v?5R�P�����]'u�����r�gp��rY��ej2��ʔ����|v�	�I�)N7���W�x��@��K�MH��m I�>ZB�!�XtP9�43�4J��G6�Su�o�aT�cר>^Q�����|�4s�����.���0-jk�p>ϕ[P�#DJW��؄_y��^��YF2H�?�C>AX3��Ѣ��L+<bZ�h�M�y�rF��x�0�(��c������T�\t�����=�U�K�QM�7 �zSQ�
�]��V������������n�ԳLU��d��1��P貞��g-�'N����ꎯ�<6\}�k
*S�٧,�ɸ��(̌g'� ����h���s ��0���:3.8w��=,^��,n��i.���l;������ǎ��k'�����XlxVHYEB    4089     e40[�q�`���f����:+����.2���%A��f��2��b�Y�t�q�+�`������(�H����,�Yw:8ѴrE�����1��ZG�9�����������/?�0]�ޝ���AYD$L��&��6����>:M�X~i|]��Ois�m���-�2S�GS��,Sj�uh��q|��E{�Պ!Xr���Ck�eP� m���t���vw��[�
+\y4]����?��S���q;y�͡���|����B`щ���5���@�y�+�l��9��`?杉B�����/W���Yժ���/b���s`������x'C=>��X�Н�4�_Z��{Qd�Ҝ+q �'P�
G�' +���I� B�ژ����e�ȹ��Ibͮ��AՉ^&eqQ��a����W/躨�|��4�fNo� �ĉ����z< �����bSG�V�v==�K�8Z�.��l�:�K��+L�< }���ϵ>h9�%�[��3(�Κ�͊��vA����L��� J�%Y���E����-��+fl��]Z�4vM;�҈Sѝ��������@�>k�@�R�����+��2���
�����`��Jj7A��%����kvJ����P�����E�83�B��%r{�^0n�i�V�Gt�� �$9�/Ӊ-5˫GV�P�}�v��0�j�c��}R]�]XB� �O����y���'��W~���rM,TjE~�1XP���?5[S��T��?)���ֆ;!��Xl��3dE���`�J�'r�?�4�����iz_;��g.3�M����� ���DY`�
�,z3�B�~ rW9/{���9m)�HTMuӷ�J�:U� ���\�����?���0�\�9��(��I9eo��nQ؍ܞ�
�������(县�5�w'"�r�?� 1 �����!���r��KP�X.R��b�)m!{���~�n@H ����h��;��������s\�}�K�JzuˮX߸ޣ�{z^E�w,�}b��첚cH6Ԩ��,16����_�׋�b�K!��K�LM���-LĐ�`�S��4��o܁ѷ)��gې~qG�,L��Q��K����i��$W˾2�+�P�����/��&Ø@8��ivi��F�CU�KX�#3��{:xS��;+��q���k����Xߙ�����C�H+��7����%�
Z�{v�2p���"���Fj���qx  �\�"R��+�pM;����hdٱgl2j�����}��sW?T��s�,!��{�`�(3�Ua���ғ{l5�Wk�)ijN?� ���#���iùz�����UζϠ��$W�}Rȝ�r��@Y�Ug����5��\B�I�q����x��s���f�r۸�<��q>�G!	�k�aE���#Jp"�~"�u���'��$��_X$�1`�_�:^C=�ݘ3���dM�)�$�#Ɗ��-�樆6�o����	���o5xK�����N�F}������`^I��O�Y�����G����D�܇������i�Q���_ G*D��pD��/����kkS���k��kю�!c�!u����R��GEh�;t�����^�\�� v���C̔"��Ik{u\�`g���\�J��VzS�c�:MfTݪ 5�er�)�2J��Q=%B���w�ؘ��R�E�F���vp�i���=� <"�U㘄a�E(�)�4�t�XO@@�(��0�ۢFb��T;�t��	�(ۯɋ/���O���F��0��ݬ�|���~������V�I�S�%�iq�+���q�HL&db���|R|�|��a�$d���r�-�st�`��5�80�A���?�T���w"��z�V�t&�B�Kf��1�Tn�U��l��n�kjks�|��nlG� �}�B\Nyܭ/?<�xήN2�4��F��e?�O�ه���M7e1��X�㽂�ë���5���j����"@��m�h,�!�k����D �QK�����{*���i�@��.A�����nyjs�#OT��p?�' ������Qݧ4F�q�­��~�B�b��u����])�o}~��a�p[��		02�]L~\�J�_�g���O[�LkOY���5��0Ŋ�ө^3�z�`5�2���)��9��-����ĳE�{x��D��ژ4Iu��������s�z����x�?^��W��X�Kʑ��j\�'�^|���O���ia9IÞP�k�/2f�ޘ-�9$ЈԤg���R�O"Ģ����I�&�����j�b'IDj��+Wߜr�)�|cv�5��R|�9��}����'rPޢ��C1*��>�E���\�����m���!�/��k˘ݧ��_[��M��_�M�0������y]ԅg<�",�����n���lCfxs�k;����s�ۼ�#�3�x�~w�����mԮ��f�f�Y�9S�k�t0����{bLb��@�����]@^����	�c7�+��v�$�a?+r�;qŷ�W	�%��C�`�p��ٸ�,fxO��]�"�pך� n"f$�����Zu:���]#1�J�Nޗ[�JqZ���t�F�� !�%ɀQ����'n6�X�x֭%��:��,3HI���qO�v��������$��-��(�h=M/���������H:�l-�=<�����n�t2@T7�D�R|��\,h�H����s��0 �z?�יlf�M-�޾f#H��扭=���)@����n}칿��K8:�-�MZ��4� �C�ѣ�:�i�����w�8L�Lq�azS�$�o?]�1�6��@�|j��2������Y5&{'�X;T"�X���͡k������K�W쪝z���7q��gwB��'�秢%��ȼǉ��M��]�!��\j���y_��a�f���pk��<Չ��ƒw�2�H�[4,�L^+��[�L^<��zwS7�u�����R#��=S��� B�I����c�#��`�g6���w�	�����!l"5���f_���C�L��M.�� dz��V^����k��Բ�q!��:����1�r�^o�V;s=WIT��� G���ҋ��~/X��[i#�(:��5e�.D��5��7�}J���m�l;�|ak�]��M���%�8����T@LG�rwwĖk��������k] ���r�~5AB3Y�sf��i}]	��[���N�!f ����2G.w+W��Xtw(
GxJ��u@J��A���j���XN����UMao�1o"�l��	��l.$�#P^X
���c(�*��ض���z�ٹH�P�:'�]O���g׸E�3��4���^�K��~े�n4d&�o����.�pT�?pT��\C֭Q��]���6�ę��Mj�N$O�í��ː�R�]���ndU���{�y����!pts(���Fd�+)b+�(3|6�ʁc��+%�.�rN�F��*ERu}kK� ԰�$��§Mfݒ�=|&!*��L3j���-���bQ����[��NʩWs1Ȝ4D�d���&
�� ��x��mhe:���q� �<��zr��F�B���3,t_