XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���rm(RR�tPO^/��f3&��q?�sR��t��j�����LY �-ERD�����|�}X�@���n�r'�zݻ�u%�k��q��.ߝ�ĥS�s����"���b6JP���h#Z�C�����$���}9S�lZ�z����8�yp;n$Ӑ\�N~����	5O�y�c���yi�����+���" �M���q|sɚs(������>`�ȏ�W�AZp1�k��c���e�a�BNk̚V�\�W+}$�n��3[$��K� l%�n�a`�4x���L���u�C��~���W}/VU�Щpް�$����V?�׀�G�MGI����;�)MNE�D��WQ�ɣ��y��t>�`FىX8�n��� ��99��Y�:���㊛�ݺ~i��H|6wa���>���_������a۸�6�ڧnD����p�`A�wc��D�RS�a���e�Q�Q���]�����=�0#�.�lh��3���I�SŚD����F��x�b/j[x���z�f�����Ă0*��]!W�`D��T�/s����]?i�*/�;��fҥ	4��Ğ`��6��DN���U���iѿ�1��ڕqChME_(�!�b�c��x˼F^Z
��IV�o�j/TNuY~,*昅���o�MYO��S���� �`����۱�re�"3��D2l�%zS��A�[�n��5�Z�bn����b�ɪ�&qt��-%��Kx��+C�Jc;t�ni���vXlxVHYEB    fa00    2260���$�!��E}Ow ;P��?�--Hy��6��s���b6����A桌x��Cv�I+�3|F6�#[� �]�[��h�k��ʐ�@ȀY��!�8��.����{>�w�!|����k�K��.�rUC��	�?��^�q%�[�ܥ�������{��N�=����vԧ�>�*�+�ʩs�����HkZ1��\l.�?�r��O
�ub����5c�����p�?���)(}����I�>�6y���� �p�p��f� �D4��K��c���U`m{��A1��fDN���l�;ꞓ+s@����ϭ?�Gh���J��]�w-�����b� �������w@%1(y��J�ku>.f�[�1��"1q���S(ή���`;�o=#3q�O�����J�r�1o{�u����]5Q#Ijo��r������fZ܃5��AT6:�3	Es	7�Kz���A��tH�)a�+Ce!�jz����=�$=G�<����r���������t�9"�<=ߞ6ׇ�Q��my���H�}f�b����z�l����I�9�ם��^�8-��d���Q���㌴�D�5ё�P1�SL%Q�[&cDvP@w��F�q��p�=#�v���o'��j �Tvco/LǪV;m�ၾ����T&��Fk��G� |�l������wJ7�SR��K]v9z�ei5�Q[UV�a�_���M~�&Ei�O�J�/*ag��:ɦ���8^'��������wXu���\�5"jry��Ѭ���XxҬ˿�����<Ӫ/w�ZY��&3kP�b��dÅ����I���;E!���K��st��e-�8��?��\x��:�,CG�m�����M� O�J�5�YG	��in	"�R�(��C����f�Z,r��%��Rc#�G��r��g����.��R;����#/�-g5j���S�8($���]_��4� �x�@.��RiBQ>(�W&�C���)�#�i��t	^up\

����o-�^y���c��_-VR��N�����9Pk��t��t�A4W #<�8{�JB�Wfv�_k��&N�h��5���l�`ΝL[��(�r���lz�ט��]�J�mS5���E)�p�&mJ�9��m:�����Q���u1V���?0q���^Cn���V�]��C���<��yR�*�W=P���� 
c��!רI��^ǡ/�`��$�A=r�.����<��N�!c%���CaYKݷmU;��'����t<��d�f�6
!CG�Ȏ���j̎j�S�� � h��s���jf���*醵��j|"�=�����Q1��A��D�����=�5�h�%����Xϧ�a\&���[i�i�h��U0���T���J���/�-����P�
[*��2a:����-�M1kj���g1��(,��'I݇��^��_u���*�.�V�A>�*�عrU���W*MĞ���ېI��r���F��`�u)��D ��$�͉8*bq�r�K��;�Ζ-wװ��y;���t^��A��0%My҅�aN3�/<3�11e�$�w�$j�=��qC��:�xhI>MBӚY��&�&c&`o{�/I	7��ηc��5%��cF�f����3�L�N؛%�����#dRI>�CMMD�zD@(e���0�+�X��Cm�����3B[PĶ��Q ]}ZuAM��M�\3D�(6�SQ�N��C�D"ђ�u�Ϥ�q�o��f��"�TǨ�d/���{-�z��aR6���N`�I��Us� '-��%� �-")�J�QҒ�ƹ|����Ѩ
�&�|��4��^|;ױ^��Y,�/��Yl���h��uH�7᢮��@��l�-d:�VB�*��~;�;	�X! ���pQԷy�F*׌�fE
�����#���|h���N�9���Ѐ6<�bI�*99m�d/'�ݎOf��>L`��^����U��u5n������`2V��t�+Y>˴
���І�V ��l!���ys�(��$-��k�^��r�T~�ڄ�zW�<��e&E�2��5����i���;e��+�)1c1*�kR.�=H�ϧ�-�+[,o��С���p��J��"��H�z�8���_���,�����q�cy����yv��4H��՗��hNy��u�p).�S	^��
M~�� ��C������ks�Y���H���B�_>�G+� �Y.��U?��X��rȶ�l�Iӝg�"��s��C^y��m��Q@�A�D�+o~�싂C�=���ku��hTF���w�@�L��D�x>,%�d��ָ�����ӱ75��cV��Wg=�_ԯ�8��\z!����[,��z� A'tw�1#9�W��$yV�`����zW��~�����L�ac�դ�2}O�V�7L�͜����&2%�,��p����C��CM+Ù����� ?�!	���i3� 
�b�=]�hxx���g�@S���g]Y4 -:Z��\>q0ڤ�Β6^G���D�;������b��#;I8����C63��&7 �+
-&*!�EN���g!��n��p��c�t�K�ʙn�=�z���<�����stn>p�.�b���.�Xvs}?�'�)f��6�J�J��"�G:0��wm�#�V�e!$1�R{�m���p"��PL
�+�S����SDI`��#-��sÅ(zyB��r��&WܗO��r�U�ј���0$<� VJj�r�hɔ�1���$�<P�`���I�필M��O�G�ǌ?RHw�H�;_�J�{�������t��n:~�L��8k�NU��T��2�u�?�Ж��ڡ7���q]�X��f�`�1,9q�Q-yM?�}�7.�b�^��\� ���33��#�@:��F|���Gv>U����&�D%s!�k�K��q$���W��s��R��� ܂��Q�*��ބK�_�s��S=R����;A%�\s|�p�f���� *�l�:f� ���G��ƒFB�>���]A?=�Ÿ�"�-O?�d@���8ח��AnA��\A�X�'�!�$>��|ݒ�ﭘĭ����n���E��c+���^�.�L��e����&.�GN3�sl"��ہQ�+a��U�w�~���޴&�J��+��sZ�ӿ:�QX[�=ݡ��p^7#il$�����
����q�F��k%p(u�{_}A,AM)p@��+j�TR�9�N��Q�M��-8��'��᫇
X��@�-\�u�v�$ ��dNbئ<�"k�\�ُ�i�E�p�?���^��9����%��!!e��/)Pv��p���P��s�S�7�^h3���hw�u���Z�
�jd��ٽ��|6ױ��V+2HE�5m���@�^�k	<9�S��B��5ݙ͒��)�M���PS�����;V�Q��}6�����˟��o:���<�\*��R.'��C���r�ڨ"g�t��_zk��B�d�J9����+e,tUq��t,�	X�R�g�-������؉-<?+*lQP��*�1]�	'�����:�{Kg񾪟M�Iq��b�9,#F�K�Mu8Ж��뇈�J���)�J�c�<}��=)4�����C�5���DkJ���z;��n[�'�D��Y*YJM�M�B�uxUT���G��6��"��}&3�K:t\ ��3��&6�����l��ߨ�yJ��e�Ϡ�C����h)/6�!�"��&�t(1\?�A0���}��2~v���NʩbձR��&W�$���v֑�E��`��~s�����L������.53S���S?x�X���r�1���~�Duc�F�������j�0LT,m�7��"!c��q���(���9�^e�f�
q9:z�6�)�G�6Hx����oSCs}�����_h`.|Ms�t����Ȋ��r��h���F9��Z����O���k�f���,�J)�[_e��w���2���ւ�iq�B�8Ԁ��B������}���N�g��i�t�ܺ��*���՞�x�������){88��AIq�o|�Bbj�o׋�t����{���-����]�����[�B����ax=�$.�ٵ\�*.X��ؿ�c=���%K����D)��+В6�g�Bo�W�}9��C�3�!���R���F*��xw؈e5g�Kfw⯉2�iԟ0�k�����D|�4 ��~��LQ[o���p���U0���> �'5�5�m�Gl_�� �>��<�F��R�������t�.��鏲��!@�C��Qt}�{�/�7;R��jP���DY���\C->���2�qP��	�֮\�m�2���9<b��lg����=P��?�������>���i�̩� JOօ<7g����5kK�n�S�U�f���9�������[t-ȇ�����F�Tu=���գ�|����3wԶ�J<�&#R钎E;��D�T�����.\�� ,1S��ʎ	ro��b���J�~�5ao5��� �z
u��q�Ȏ|�M�B�'"�[��V��(<�(��h祐u���h�#�{���E8p`��Gh�J��9C�h�Lm�m�)�=����dlr���:[�H�����j�O��U;o��尙W���h�	��W��iA?�̨�4�!>�S	W)x�j"��dx��W\����h�ݫ�_	�B�G����?��}\3�-
��Zx6�Y:U�^48� f�c;[��w��d'f�C?&@�Hm=�S�����Ǿ?ye�O��,��<®���̲#��KW:��R1oV����<��d�#�j���ƣ9� ��v|��B�Jv�b������f�%�\����vE�� �@�����c�a�1��y��pNWT�^����c��^hh�`C��}$�Ļ%� �7�t��mu/�j[�J��-�:M��b��^>�����b� F�0B���?�=8r
=���s
*��#�D�6?BF�J<���M�	Re�@���쑳���zrg	>�W�;>R������_���*I��(0��`�<�R(�".9��E9	���L�X��tT�A������Ý�|	��&`��}����n���{sk5���	�)����4�����7�� � �b���p.|���&�d����m�cC6�|i/A��Y6+!2Ԡ�F��^�kʸ�����B=ȭ���K��a��r]<�<K�΢�W�ђF3�a�>����L��n`��/�~P�V�Z���2%.k�̅t\<U3Nu�J����	t��*��i�{I���������Y;�����	����(4n��_~�Zڢ�'�vo�//"]r	�,���� Kq1�%������A�U7^��'�^:���?F��`���H�Y�ǅl)I?E��H����@�I���Y�UH}��A�?1��	ߤ�'
v�Y����z��@ԴT�0R�ہ��[	��i���zJ*_�(�J������w��b�9]kS��'Ϻ9�Y��,���G��lq2��Nܯ�I�]��|-������6�!�Ұ������R,DOd�[V�k�$�/N� ��vzͪ�on����nJŐ���N�RnȦ��VD<ԕ�=׷�K��"ʴ�LΠ��aݜP�����__�M\�����{0psLi�����b���Z=}:�DO�W�B8XB����O`ٞU��#�l]��+��q����o���T�`�Gd�8D�{i�7;����A��ݳ��L܁�s/����bG��3ъ�v��
����o$�317Z���	S���Ut��%-t����ȳ$m/���{�)f�Ɍ��;���;?��#0��@�q������Й�ҋ�6�G`�Y*���b�h�ȑ ��p2�V�eO��y5��k�5��$���>����,�H68��mA�V�F���3��C�-�kc�#7N�.g�\�q����]� �/{�RXX��j(�$٧
��}��b��l�j}�$<�f��n���~�R1��xԣ��%���&�T��vb�n<�� ���}Z��'$+���+���bs ��GT�� �K�rNiZ��D-���zz�`bڗ.?ӡ�����~pX勩g�(�ͩ|����v,9\�먜V�U�~0�9	<�2�˝�S�(ʊ�A[ӫ-�/��k��������pzhoU��`$�7xqe�O+$q�r;s��»�e2=
9��tu�l�W�5j��
ʪ9�d�͐�f`I)��j��t�� �Q�����U3�i2gE>�"�$I�����e���~.�m���V�N�����1��*9Cz0L�̀�4k��$���x�eӱ0�PE�4����j�,�}�eG�!�SWI_2����vdu���:C�T���`��.;P8ū6��b���2δ2�7�G嚖�=����3mr�nM�*!�@��h�##gUK�7���ڷ���~�ܪ�FRq��{�'G*ޤ�{@(R_�;wS'�f�.�
 p�~�Q1�����U�h����o}U^��
�.�}@��!*l	�M����W�R=�7amr��g�p��%�^\U_,�(?hJ����~���8R_�N��+�:Ve���=�Z�t��jۋy����+@ʏmd:M١XAN;U��(�kP��y:3 e�*��?!y|& ���	И�+�	����b\�Ԃ]�k�6E�g���b��{���\����r�Rt$�Z���`���A���F�8b�j��D�^{`������������z|���@��q��已���>��#2�!+�[hR$g�O�=���Y�E����h��<%����r��![�yh#O7"�	�}`�w)�/���*	'4�����k?�oa�.򶛚cs�M��o?e9�, [D/��gjcY9�%g�~z�O�;GCk��CN�c�8�֮�'�g9�_�)Z��â�NBT�с���hsSԙ��a�� ��c>���s�@9g���(�B�9�ÐT~����)x�@�u��'"�W��O��O�/s;��/��mh�??�Z������3d�J298[��P�PH1�[���[	}��9�Y|)��L������-�0��.����>�{yԭ�N����F>������WL�E���N��m�	����o�q�f�����9�|?� #f�R��c�����
%ç#M[q]'x�ֆ>�D,i,��({J��]���X�(�@J��O?���B��j�aY�1�ۼ�\�t�/�#���D�m���0i}����1[i�SIzF�D���1_����UuM5F���_I�DO�Vkz��-I'��z��E-�2=�]�Jq��iI�0���xFL)���1+东wgC�Y���U<���D�,"VS�P؉=Z`D�.0IU�ժ������'����Ơ{�)��%w����#%:����p`8���#3#���@���۽P��,�~��I��VF���3�e��"�2D����ۦ:�����q���T�����g�*VK��W$Ղȝ1�w�����j�,��1�����?�
+W�(��9K�05��9 �Q��2�p;hf���ўWL���>��o0V���^�]d&�Ŧ�Dl ;/a(�.�}�K#�J��]�r^^Yɟ��}�8l��P�I��"���@s1�O/��p�'�FZ�dt�p�uH� �*vK'2�%�y_k,�=Tj�C.f��$*��7�q�͗koq�Y��$;�^�����T턢 >��CQ05�,�uh��`k"��9y�� L��|�O���Ds��ڹ�O��K�ڧ�J�miO~0���Y��j�ǝY��m|�ËY���8�D0�Bm�t��fu����9��6��tb����@����W�)�q��ks�	5/��^��A��p\�J~�d���k�8C���'X����#���I۟=��30����Y �Z΄}�>_��N�YY,��v/ ]�@��w�ѯTnw��V1η�ku�=�j�p�� v����!��LL4��#��8K���`�{rl�b�M�aّr�8�֤i�K�E<z���p÷��aW���x�o0��c�7��g�G��tjW�B�ݶ�����r�]%I��9d��*Q�u�	���%J�H+Ӹ����å|3�_�넺��=ƌ�
hm,:ӭ�M��/9���M�%n8��� � �6���F��^?(O3�>��rMn�TE��_�&�Thcj�=" (N��h7 c����xI�-�����8�F��ZD����ې���}����;$"	���jR<:	��<�c���r]���z�ƫ�R�d҃QV0���!X)���e�3�NUaDK}ә|@����N��>Ɨ_��
,4��ʚ�v�I=�~e;���WD�#����$�y(����M��Vת���c{Hڷ������h-�G�@f���k%OH�q �8U��,�ɕ��2�&1R۵"�:Q~���/�wq�jJ{ߗg����B&`��K����7c��V�!t����?4Q��K�K�ߵ(l�~l��s��M�WJ�s�xT��Ql�(��`��]�F��K
�(�I�2�eU>��|�T��K}���eq��J��(y�>t�n}��%NV?����(TMq�����3�ql�܉���167���p?	
�(�#D�X ;�န'+L��ZI��f�N]h�g⋺� +g>H_�½�����Ԧ���)XlxVHYEB    674c     5c0F��J��H��VsϺ���
@�G�+#�UJ��z��j��*����L� �c�G��Q� I"{���]�h����������}��y�Cֵ��T�tnz�8�0���}$8ي���Z[���SU:!c�/+J�x���F�FOJ����w�rq"�^ ��DW7�EC�#����yO'�[���K��O�&�_ q&2d�gP.v~��qS���\��P�� {�р
kE�5k���,D$a�$�)����C{��ڎ=���O�y��N��P1����j{Z3O�K�(h$P�e[�W��"V�?ٗnW(:7��H���� ԢI�J����Z�a�Q��*4���͗�/`sEɋ���}D�C5r}��NhX���5��H�Qz�E�6;0u�$~�v�'�R��<'̋��+�K�0��A�7
�Ky�^{~D2.���N�W�$ �y� �DLU�K���WIO°�a����Z)��ͤ���5��r��M̵���)OR��f�#e^� 5���ko6�CoRu3ź~��U��D?����h�З���)8E����=mU�H7��dh���l�ɄT��P�ty]��g9HHAF�V�dv�ԕp	�V5�nB�T�rB܋��*��/�㯾��=>�M�N[	�Ȯ��φ�PY���6�qzГZ%ў"X�v�dO�Ӹ�B<;[i��qm5SKw@��=�$'H��(�"���z}�\�Gե�;���5%ZǨ=o��F^O������p�[]-��Z!��ϡ��	V����]#v�:"�p VA6W��@�F�F�Jzuh��!f��qqL��p�3��"���uRx�Z ���^x�'��m+f�L@���r����F� �h5��i�>�V�O?��@Ɓf'��P�n���7��cR-��aU�\����R��s�ֈ�S�N�f��N%0.]W� ��~!��@�`���W����8R@>�(8����G����|b\��]���Y߳P��Ǫ�?q��9�FƟ|`�q.'��m�A��NyO0kr���d��r�>q�C9Ћ�X9���h};�p���:H�b�lf�;��9�oV\5�F�|�a��b�
Q��ZĻ'��U�d]���q����j��3�O`�B"��S2�~��W�	H�K�"ǣ�����ţ	�P,�^��B4�
0�}'��s*�tRP1`,�t�/�"A{N�����U~�����wꥥ(�ا��V�/�3�{v��	#$�I�m]���k�C�C�@܋��2c��d��+`�~�Ҟ�L}�R�b�m��,f5{W�\,EE ���ҒwI�	�\�eD�u;>��0_D�P�S�mM�ۙ����� #@31M;��!�5o0�T&����
��,H��-�F�NrX���F�ױ�I�!�l���zO�E�0ɚ��[>r]���l5���٢����}�w6�ɷ�9: