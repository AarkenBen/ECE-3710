XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����*_�5&6(Y�#���t�$}R�VrT��)�"�̤�#絇�9H��z'���W)�V���i�N��:����B��0_�>Dc9�1����̰@A�c���Ū�7,x��'*S���IbH�A'�VPgl�_{��,-b�J�HM��V�۞h�h���Z��{I�4wmMu���#��ܹY��b�Ƒ~���3u���;m"L�5bX�������a�����кp�(����m� �ص��e�pK��A8�<�v��Y��o�y��`��v�m^r���S�L��?'ͮD0�~�������C�R��<]������ǐ2'���qՌriG����Ǜp4.W	��K:�ʍm�2���`��Wo�yF�Ve�v��>In	���ßm/��H�va�(kdtZ:���s
����b|0�g|�����]��N��@�y%�ܹ��}���Ip@�>�ӐZ�h=�+^���h���Ud�e؉��'ǔ,��6��)-�5�0�ot���VR�� ���혙�UW57�9b��&em��ߑ%N��Q+���S^4nV��>���{5�UKے����FPN���� 5A֫`S)1��݃΍F��v��\��\Ĭ������x�dZ���_k��1@�V<��IMm�x�*���h�/qP1ce`�7�9Ù*Y,�;75w���/�����5��p�
@��63������=�۽4��j�V%)�g�Jܲ�	�P�ͺyWv,���a��[XlxVHYEB    9de1    1670����V]�����9j�R5��#�ĨKޜ���g:z1�X���<��w��~�����C��G9���F��y������L��R�p��X�|a]0� ��eN��n5�I�rPE��o�ޮ��?x��u����@5 �l;�'��;B;��)t��tG�	���ޒ3�Q5JIx�C0~#�i��%7��߹u?g�i�WIru!n��F�`����[
:A��<�s��͌`��K��RT[);����)b�x�u�)1!X~5b�bQr~�v��z��h.���V5�X��i1G]�dX��T5�%�A/w>��Y��ʈ�r	])]�5r�sl�A�ta �&>ŗ�#��N�F�⶘����eHv�\ͼM���s"⃦�Y�P�
�|].۞�n�Je%m�@UO��nb�҆s=�Ǉ�Ys<���3���p�d��#��yf�����c��I��r��&�6�Ǿx�P�H!L����Dh��K`�tX3�ؚdK�_��*tv>%b�L�qA��Y,��'��oy��zj�	�7#��k"F���?&g�u�#gˮA���k�z�I�T��0$7!F��6�A�>�EVϽ"IB_��oZ��mծ�-�6@��y;��d��Be�v��<#C�w{N� �B�l9���	��'��J�I+d�\����T2A�M�ņ$�qOVe�=�QU�0�|aO���7^lj��n7vL˰�x��^�W+��`�\� `Ui�U�Q�� =t!gm�Ԭ7�]L�T��FD:��#8�Ga��c�"��X���<A1aX��a\����q]��>-6�9Dkm�=�A��a�,nG��� !�c�0֛�.�.�^Q]ɈVy(#�x޴�SuuAAd�A-ܵO�T�n�x�k�W�T�>Tr��^�Ur+��2���Y�	c+���O�)>0�	�@>����si�X���B�o��>PƳ*���9+�K�"K�i�E��ꖜ\��[x����(�
0!d��R�3� pR�BCG����C���(�N0OKW�A�4�t�y�o4n
�AG)�aCh�w����V�l���H �h$�=�{����c������B}�>x�����)�,X�ҽce�����%8�S��
)E��G���)�Hv����#�
�����Y��]$"!��7 Lmu�01�/-ků<f0�q�Mv�r>����5�T�Z�]��0N�VŸM�������q{��	˳2��-~?� �2:�����GE�]��H������'���&iq�S��}�y�Tp�S��x�f-k�'��;4�~���t&Oۍ�Q��%���
�~�ơH�>\z1iz��a|�󤖴��P��R��}ƽ˸[5��9���A�,���	��N��ĺ$g���>�H����1�}�B^���gkK��_ܙy1@#Io���2�U��H��rH�P�2]��4��"蜳L`�Q�I��8y�����e&4�M���	]Az/B��G�O��%�cp쯪Wb(��v�W�1�9 �!bP��z�IS��s&}�o�$!L��5��.�6�<��E�ip�(�
���� BH�]f��T�p��CQ4>�j{�K��r��pU�J�."�-�/�{�߱G>C�N�2�M@MS��h&�/M�G[�?ۃ+Z9y��b���$)����$)7b_���)�Wg��S��k/?�gDۯp���1����6C�?��:o��ƌ�̳�^^�Npo�c:�\9���B~b)���	,6��(G.�3f��
|S��`��VG����<%�Ã��YA��s��8�W�AWq5V��/�z}8��w��a1�~ۊ�Q���H5z̋����^>*�%BƬ��P��;P-��N`1��N�;���P�53>�a���MX\S����j.O����a;4�G��yꗹ쁂��kewbTT��+g2ᙓ�BC�o=&O���{1s��f`o��\��c��0���ͷ%-��H���xǲ��/j�vc�� �<�XE�^�~�ǙƎ������qP�f`�O�v4SڰP�ܵ��:	h�sH�U�E�:��'�&kC�ˎ
��~%��j�T,�s��o�Gq �i�Uܢ��+ݎ��o�R�2=�����ۿ�1��e|I��V���VU�)-���\pk�� ��m�qDeYCN<i��'���_x\t����8E�'�����(xw���o4Acj����`�N�2��G
-u��\*Ǚl*���>j�#c�yϡ�.��WL\�Nݣsm����b)0ckZć���C9�q#���!�tq�Y�|������k����͑�^��[ꈟ��R��#;m�[��X�'`j>J0��\�Ʋ�M�	���&�		�b��y�5_�Zfw8bДF0L�b$�;"w�Q"����]3�ƥ���>�V]А��Ӎ�{9��tO��4%]E��`�
4-V5���%}c+ ����F�TlI���R�Bt0��q�1F>2�B�A�2a����'��"���W7�T����Ow�7����.t�M��=�^޷a��[�IL$'���7��.Fm'5�m�۽s��I�;�@�1��?H\�#ˬ3�e�|f�c�`�`��f�27)!�7y����������t�r�#T�����]t�	l����C�tP�&	x:�U�\ݞ�(R�~�Pc���J�|@�5MԳh|Մ��b�C�ҝ�E2H��|Pµ��;f��m�H��ss�/�L'����z��bΞ�����
�$hKf�:2�Pp�Z�1��Y�=��{��s�Jiz9��l�˒��,���p�Jv��F%���l�_ @��e�tkI#�wUT��������n�@��<��^�
�����z ��&�9���^�b �����e(X��2�e�#ÿz{�dQS��7:8�'r��;�\�*��H)�+��u_�͆��هo��]�v����W���!����t���zƍ����=I��#h��g���Wm(K�w�,��[�Lp&E�/8�wj�V5�.�|[�7�>��$��}o�t��9,�w����Z#��Ӓ4.s&Vv���|r���B��jBU�a2�ĉ��W�5��h+��ň8��E��GJ�V��Z�w'4����n�.c�k޽h�o�hv&F�>��	�"��y�_��P� 51���+�;�t��o�T9�)����[/9j�h¸��{�vb������	ɣUφH�E�B�����д���{so6�,��ų���p�����ϡ�����ia׽[J�,�$����*a�Y�����G��0��܁��?s�i�}_��֝Y��z�Q2(W�<�f�y�[�����m�*��;O\*ƋG����`��N'�쀎4l�"U���ނk��KD�5q�C�f�f����B���u!gg,�j5rU��zy���BS�� �ƫB�Z�C��7̻��	��n��Tf��R��т@��<f���!pb�^|;���{~��u��T!'��0c>����4��y 
�]/�aBK����-���{���iq��������Vwº��~?�h��Ǥ�ZǓ�;,���-����*t��%�N�ﾭdX�=|'�v#�q:�K;w���C�c��7� Y������d�NC�Q��h��}������>@�]r��"a��S��ƹ2�"��OF:ɨ����0�=N���U� e�j�pVZ�s�חk2DX�U��@=��9b��{�����Ҋ�{Zo����@.�9���-1���3��)�:6v�Cf�E��Y�,�ѳ6Dt�n4�Y�>��!��i�V����1����t$�q2O*�Z�<��4����n1l��#&�3����I�j�����H�T�[V�1L^��D8�����1��������剉9�w��{;���e�Any��Mo�^�T_n�2�5���k�o�	�@*뫼R0�-�ki�2݂۸^*gx]�`�U&�2�m�����*%�LO Y�-�r�Rw�Xb�6*(��V͛�s�c����o��r�h����g�ݐ(톉��9;�Tg�e_ҒJ�jj�{n�b�� ��D�=�^���)�{�0�Q�t��a1>��f�`����k����țhGţ�I*��vE{}y�;�׫�39��8���!�t���iDt�T�w(���#y�$T*-\�^�3���+�fP���^�|�I*C#��s/"5�3�Y�XE1M����j�T��B
��g):�T 蒟cPZ����>��d�7	G�� :��L,�C�A�y�MaO��t���n+%�ÉP�Sbp����ܦ��T,�a�pZ[qT1�i\a�u_�&��	V�{�&23�%����.P�#i�T�S��M�X�e-N\�a���t5L^�q4]f��tY��qk����ra�3�����P�g��^hj���"i��Sw#��UȪ�E�3쒮{�c�:�B�����~���f��,��LO�cM�4S���w�Sl�B������Q�c*��}j�v8
�%�n����T���}V*R�c!-�q�����.��1*�8d�+�P6T��<$��798kx�&&3Z�\{Gji�%��@m*��:�$�C�T���ƆS�&S&�U�>��m��?���4؏�3�Cż,u���w��0j��N�F��AN��9k�Uam`������@���׽�ٽ�g֛�1�
R=(n��)��Qy������DQڀq~�P��]d@Huq۳�f�G�������\H�|U�Ŋ���Oى��	R2����h̜�|f��B����_�n��rV��2�+/�J��bZ���\��J���Ѐ�B�/���>��=�^��Tl�:WU1$��5���8����3�������[��7w�"j���M�miy]
�˹ֱ��5�"{%;�	���8(	'�[z��f�4ݢ�t<8�Gs����h�4cҪ0zN�A��d~Z��t �� �nYQV�(vg�r�P��5��:|F��Q�-bH|�+qOR�㜽�pX�T���x����������r����I�(��jn���"e�����w�t���ʏ�2�R�D5iNXa��c+��
W���Z_c9~��½B9�n՘��l�Í�?Ҡ�����A����\�)�WzԱ��LŠ�I�d\�?�->������o*���T��G^���Icf���Rc�WW�p4w/�ء�]1#-���ٸ�J�U+����V1%F�����=�4�P���p5��
�������=�5d��H=��WR#C@k�%[�����]xz���{陀�r��'-4;���Mc�4f�����h�C�B[
$\����NM0�4�R����M��o/~C�p"b��=�Z��-b	�-����7J�B����A�y�rGR��m*<}��g!.���!�Z�5:Z�f���ɻ���_P�ǝڝ��ˇ�D��
�]_;50�`��j w�u�9'-µ"�;P�@�a�#���{?/�*�$�F��Y���p�!�Ǳ-�_�<uB�X����@��5�5��,	 0,�J$��׮a?;*�p2�s7�.`�!	~��WP��/�����8�sϵ�៍�L��+m�-�Hd9��p�+)�Z0N.:[[t\D_]�5Ãa�׷� �wB�]%fe�u��G*;�s�隁+�BUe�