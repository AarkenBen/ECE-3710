XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;j5�DwZ��{6�����gs/=�/%	�y5j��l-��1pWwݙ�+!qU�g�Lf�iJ�{�s��)�
��-)�掳vg���#�����b���L��O@h�ɛ9^e7��r�Ξ�g/k�-@c��RXpz�L�n�3��&��֝����ob��y�}�i�|	�l�4*5�L2��cjؠ#��X�HL2�ʯ�L��S� &P_|�%=��Y����/�_��)��+�E��*�,B� � ڼ6ߩ�+0X?:f���"d�B+'�?�\���bG�tX*u12`%�M����O��I�C ���P���uI	'��1t�}��kqE�Ks-����j�`�j��{����Ym�k��  V��>"��Y�E��=�&>�0� =�Њp�ץ0ݽFyp,N����\��j>]ï �5N?��>�4W������Q�$��U�]��O`���0�X�n�X��Q��5j���|E�.#	.{��.,I��k�4nGjnO���ԚJn=��I�=�#f7����=��'vt�(�Ex�L�0#���K� �E	J�����!W�>�
�q�܌����?����������Ùv�p1��~<3T��v�	j�����9�`?�ڞNc"�-��;6��F�(������e�Si�1?�ZOi���ˌ��n�� c`UGƂA��ă��~����������1,/� Y��U�����
�� �e*�@C�\�"�O&��%�7�/�%O���$Ɉcֽ	۪XlxVHYEB    56d2    12a0'Z�0xF�f#151@&�L[��+.���⇚S���k�MW�3Yk_p�c���A�?�"n��y�%����iM0o#
�TΠ�#ut�F_8���X�P���Xxz�/��H�=u�Z¯Y�M�K�a��֫)����A̚�	�J�>Dm�ˌ��o������ŉݟC�W;b[odJ�Z�R��@���W��k����o)Z�����^."�z�DQ֓3�I��I��v�����j���m@r�� q���=t ��2��	�8}�Y>�e�?{Ve�U_�7�Nt���1���D)�93H�bOB�>���	��!ޜ��ML��ax&��P�"�)�?Ar�~����vѬ]��u�΁n���2���m��������6T8�C�\��N	�~b���,��u��II"!B9��0瘖Y�����sC���$���c=|���N�+�E�y�G#�'%"��s7�'*?�v���宗<�"�؃���v�<R��Pfg���	��LZo�`��6r�����|�.�U�ޗ7'�S�P2u�� (�wR�̗�����s�)j��Ԏ��e羆� :�܆����o:�SY<��7��{D6C�D��<�k�	"�K\�8���1Y��(<;�cN���c����w[4��.�͏v�I�j�� ���F�h�8�<%�p��G��n�W[&�0q���®�]��mZx�9�޳�����XU�����k�@�����m�^��E���;���9�����qM+6����V�h����$,��"J��B�ξ��@����#����GE]�纠��k��1�>�c��M@<�7X̰�QçWg� ���=�ZÆP�b��B�Hx��#��Z�P5�u�'�V�ܚ�e�����ъ�%t�{Љs�	�<���tmG@i(]R�H�~�؋+�*�R<�T� A�>Z��\*?@Tk�2n�(�#�L�k�$*�-2��?-��3r�����3��
����r��:����(9�v���n���#Vv�6l� /!CBi�|_�2�D�7�YЅ��v�+>ے#��!�$�;)����]�b�6Ⱥid-ȿs��+�$*q� ��O�_�� L�=,����H�o��q���[�l��5*`�d��+C}���sWx�|���)0�P,�����^[���C��V�1ud� ,Ox��K��?P|��RS&W3�S�M�c/{'�"����\Tǡ���\:���W6|ctvz���e��"���g�Xҍ��_���R�0��~B��m&8j���D���JfKTوΞHv�.��/-ӏ�Mߣ���ۯt���<~j==Ȳ2.��T7bc~{D��?q��Vz �_�����oڑz���GD�=^����m���cUF���M����\B���z)�C�M�O�X՜����I�v=a+�m>y��iĔ���L{�l��!�]�T�C,�w���e���6"�)��n�O�\��� �6a&D;dʟ6.�ږ��F|1naRKNh[���^��;�Q�kF�W�p��1z��0���Y������q�4Ә��,�>r��v[��2��M��&k��*ߩ6���{4(��f�a��V[sP���f�
ݦD�7��UVq��&	_��ɺ-�%2�������1�@hv�nW�R�D��?7eM�K�J2�T����焆�?�v�3봁}}�T|���<s���G�d!��阪�S���Sȗje�~�Xf�Р�S�v,��m!�u�p�[F��}_BdcG��<�U{���9�T�d� ����ټ�Q��e����ɀ�8q�|GY��>!�����<;���g��|`ҔE0�y��c��4̶�	���w`'~���������B:��6�մ��^c��[sr��r�8� ���X�
���U����T6+���oH~�	B���,u�[ke/1O��Je�A�.��M�^vf�=&��?�!�ц2*i��~�H>��[��i�U�`�tqٗ�U��]�9;�C��/V	)��Q�ܚ��
d�ɞ)�L�M��곸��v��):��Db��/�a�B��h��T�I$H�t�:��W}�5��2�������UX��������zܒDZ	Ō�n���m��V��P��D��~0ռ��� F�g���t�2V�٤�惰C|2NP�C��+Bʻ�8�a����S�Q-�w|�>bF�uZ�~�� J����2�Q���gr)H�'��x���\*�gF=��c��>̈́@|ySd�D�؄� ]LXW�#m�"�_�����<�#>��e�u���ts�U�Zl�����ڈ��/��+e���܄�ؚ���w�ƈ��N3J�V�!5�Ǧ�t���c�cͪ%��Fy>}V�����~5|X��M<�4�NJ��񟌯�Y��%z���n�.85�Hfj��9��H��9�ykt��t�G�Ōn+,>��*�v��P���k�n!oM;����E�Х�9zXz9���eҶj�� f�[����v��s�������e�r��A'88!&��w�7�as	k̄�z�>��9����P�*��@�|����V �e*�A��(����M�z�B���_d�h׿�㛺����~0l���l$�[1
~��2��!��S��"�>h?	B����Pl��v�%K�1��E߅eO�"�����q�P��ي&A�����@z�_�1n���=cЂ�������[�o�v�K�ٔ)ӌg��X����t�M����ڔZ�����y�R��V��䕚�F�-E�\���+Z��%��'�f� Ȩ�D�Lڽ��T�d��a~��~_��逼7�<��'�k@���S?�Ν}�.���'��r����+zZn����H���fOݪ_�Vh�����R<�g(d����t'ǛB�j�r���	@ Gfs�V�k(@x,��iB7�O��*��<v8o��\�SX���x�h��Db�ʌ��h�X�h9��'r�����b'Q>����	w��ph�^���&as	�_����6���V 8ŗ{R{]�(�XgOB�»y�T1�r�݋'1��a������i�v:R�ŭD ��*��v��o�_�'�-�e�Z�����Zl���ͪ�k�C���<F3a��4�C����c�N;���}*���۪o�����4���-|AӤH���M��y����o2��u����8��7+s�"��(�<�1~���i2��AR���l��~S���4���;��#Q��G3a���!�{JJ�f���.D�����u!�����$xi�B�J�[P�q�ӫ�v���!~1�$<G/	[CSwŜ�Q.�����T��n���%Ι�n��|�ps(�$�Oa��:D�
KS(O�j.ϔ�_(�_���5��Ju�M@���������ڣ���.D06��|�2�q�՚բcڜ+o��|�B�3��g#X��˻/��6�����kD(Z�~\�q�?[��� |����[v�86��}g{]��=�>��}cO�����c��i�y���>J�Z��k=���2)g�\v{��"��2��@nl�1��<�]p*N�a.��a�Gl��h�E�T�qY�f���O��'�.��'%��M�B\5����vṑ��$*�A�����'y��֕�<"qP�Y	�}�7b�)��.��g`]�8�I�h��W8u��h�0| ����V���v]o�>��!tS^� ��\�,b��hs%��/��b���wtM
8[����MLC�q�����Nlj������q`�e��T�kܖ��ߊӑ�Z���t���"�~u�}��,t�E�[�~�h��H�i��E���t���i,�g���MwҎ�S
F���*���O�2%����HFU�lBVTX��Iǋ<�g��P��Cާ�j�J(���!>�M0����(1�#pl	jo�x?gk˽�6��A\	�gξ��mmd� �Ymp�K���3n�̵���ϛa_N���9���B����IU���2!��v!��[�� T��y���Ezs�
�z�E 	e���2������������n�ȫX�G��]�����2��U�"+�+ʚ;�4{��O_[oܳ|���"sTl��cs���i�z�yJ��Z�) �sI��/�}���
��g�#6��ub(k�n$z�oFg�t/>7\*& b�w��hI�h�������5.�a��	����IB��[2��[R
�����Վ5t@I�~²���j rGܑ�m�o�zS�r�!�/���NpPP=ڐ�cD�L�Xc���X�H�t����N�-���*@�e�ޓ<:<���	��h+B�I���K���귛�G	#8EH�4�q��p1���~s;N*J�C��w�Hh~c����w��+�B���j�:�t\w��<����Dh�jS��G�j�=�?������o�(f����sT�@5��D��)ug����i)Ϸ7�}8��ew�ǿ��4wCL����;k���G�)լ�u�4/�մQ,��^;�z��#�a$�^/��+��Eʙ�*4���D>N�3��0��T���p����z����`:7���o�"M���͏5r��� ��<�9�<(m u���˰�4u�&�@��+�,}��
��j`YLF|�W��0go��|����݄�]�!P