XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ӿ6���[�R�A� i��iz�)����(��$����h	u���B,0;���`����\c=�f�4�wà�	٥n��+��/AݳS���}��[��Vǃ�/k�}P��'�G��N�{���`>��s~\���	�}B��Z�./�G�������P�B"شK�'��w'����h�kh(*��8�S�cL�y	 �w�ݏL�N#nA��c]7@� :����}zǭ��4�#n=�! ��(�7S�v9���43��X�LOr��|u�p�%v����)�$��-����HE.���cu! ��"��?�tՠ�[���S5�j� rF����e�?D+a�G��/�
���o�6t�X6jR�5�j_ٌ i�b,Y#��W��;���c�*ytá2�,�S{ϝ�N�������~���L����π�����v@&X4:(�]1��m�lē���6��z��x۟ �E�_�.����C�� v��>*��bwX���Oe�y�7��c�D9����)��iUU��
'�<Dhz� �d:���^C}v:�P?Y����1D�׊Ns
)j	Tqn~yR�<s��p��|v�P���j�q�{]r���6�!�r��5xk�*��+�c�T��	�S�b�4�_!�l%l���f�A�cx.<DP��k���uv�����G౴�o�,�����l +��$�M
��v��g�;#d|ge���˻�H%$���5n0r�3�Mq�Ծ�����\x�|�%�XlxVHYEB    fa00    1950^��BDva&B%�nYr}�2��7[����#�t]�Ռ���!������+�@���"�*W��������B��9Fm��2U��$1���;RE'n���:��"�~���a�./3&i~�w�7t�h�%��{X�O4z(J���hP�/fr�)'1Z���* ]�	WW�|,lV.��JW�(ꊋA�_���Ϲ5����3 	�lԷ9���Z>�+�PseG� �f<nLC΁�o�?<�!�
 ��:�^�y��qr��/�}�4n g��V����D�gϑ��x{�U���<�.���k��X�Nz ��t���o��LڀDb&�U���`��9�kh��s�x��
�~��pƽ���Rn�bu� y�����"--��y��ί�-"���qQ�A�Π"DQ����cɆz~V�"�w XlZ�|��?*�p;�ޱM�n.f����qI�w���+Z���6��ԇ��?6�J?�q�� a�k�稬��֠VkIћ�����1��6aجD"���b6�M�A��)$���B^ ��\���/��׾8��sgW��˅�5;In@%s}1 ׫;����ʣc������-�ԏOl+ݎ6z�0�ڹ��I�v���pg�{�V@i
Jc�J�qB�Z�,4c%byܨ;9E��}��*�f�ˊ)�/WL= >�nm�+Gb-
S(q<��yg�~�l��	�P�TY�#�!����ě,�JR|i���c�_��ބzxs.���o��N0{�x����]��7�\X9��8���2>h(mX\_�Li	=��,IH�ٸ��� ��;-8V�"4������i��O�% ����ط�I�x<B�'L�����;"2]���G3@�&2|��,�k,�E��XϿ��	�>��7�d��XXB4��Ƶt�J8���ho�:|�3�c Wڕ/me����X���Hv܆zr��/��"�j���L�h�C�	w!�gE�Ϛ6u���&C$�����C�h`�β������
aT�q��t\A��e�Kn׭�Ȍ���n]3��\*��B����w��(����ّ�(�i�f�u�>�-�2,z��Y��;/���Yj��T�&�V�TdFWs����aCͨHH�������(����]�&ʳ�[�^�9şu����Upg�-Ks����� �9�!�&�3cۚ`��۹N�x�&*(��҄m�U�t�!��
U)2&A�2��>F�m*�e��������J��f����	���<��t�Ϫ�?�=��ݚ�C��|D`KY'�,���g�B�͝���?.ڧ�ƅ
 i��'Y�9�X�]���P�T�����N�'�ܳ�;�yvil]�Õ��-4.޵�;���/`Q7�p��'kpr����s��H'T��r�l�ڙo��!����SW')F���@T��e�0��_����u�|iGU4���4����:Ef��y�1��%�u4a�7̜Z�z�������|���|�������Q+z��3xv�!��y�י�o���k��n(���8*E.�&��9��`�d��i3D�dI=IW�dH6����h�C�2�U۩��H>^.VH�*��˵���~)�"۠���ByM?��A���r�Ԍ�����Ǡ3�~�Oa�3)E��'�9�"��YTy���a)���O��_�DUrMt����mHZJ�����AVV����OI��~��H��2� +�rgu����ܥ�x~4>�@I�>���������P��m�]�0���R @&��)��x�2�)\�{���ͨ4J���Y��������N,j9KN����E�d�&@iQ�P�Ddh�e�1��'ؙ(�ة*��n�͘�^ýtX,��R�����fSQ�,6h5��F���Q����Q[��Z,SW�['�Ɨ�s֟�X�dX'QǔR'$�=�W����8�蝤��\��O���#�!U>��|(*|f�u6�Z�K�<A�D�v7j].V��3*8L>�ؒ�<p��g�@�	���Lt���r�wb0���ž�E�5�T��:��4��w"d�}���oE)MoG�I��E���.j� �p��J.�yJ]��?�=�'�����NQ� ���]��ص�4���k�)[\�y��E��Ȕ�4�n��iYG`�i+"aݱʣ�9��-��°�@^qcDU�p�qX�98;ط�:�Re��C����F|������v!10.X������s4����'�Q�(L��g�֩����{)8GThHP���.�.������_�3s^֬�O�48#ݒ��Θv��Ĺ���ZP�}�ᱷ��2�� �0�2��qU	��c�&z�)Pr����m���A�Q�\�2��� �d-��-L}�a�q�<o��7|q�
:4۬���]�ĳ",��x�N��w�I/�[�#����=�
�"˕cf蝤.�	����n�:y�Ȱ��%;+p��� y�UN��̽�2�~7����H�,(�aTD�:kR�n�Y+J
X�����ޙ�'�����y�T�z�2��S�{�=�zM�fN�ْD�����,�A�7�)�jȧ^���gׂ#�%Ac-.oj�%%Q��dQ�Gk�^MfE􃀂�X.�n�^�ESߥuV_��i�W9z�$=��njo?\-��'�
R�.I҇�;������\4b�C�=x����;k6*���N���2;�_�X����ff3�ԇ����Ȝ-�{���E��z�6��Ӫ|vo�d5``^������� i=c�hЍ��q�?�<QW�	��3�'��p2�D�ȯЫa��.1�sѬpsD�/J�J�O�t�>0co��v�R~�/D��Z����ײ�w�	/ |�=���-T�W=/'�Nn=��FjX�7�'3W��:F��>���t�����C��D�1s8C�wXo�l���L�:���v��e�BV��9��3!m>S2�f[( (���-�8���ި��Nj�#��K�@BSD�ɬ1!y�k�)Z=����r�l��ŧ����7e����6p��g����3.ʚ4zb��ք����.F�J���f��}n�̰/��$�F"p q�8����)�(Յ.�qtV��!�-�pV%Q�1Q��j<�^E�Z�1�q2@��ڹ3|~��FT�ց[\�������e���e�9!�=���؍�`T�6b6�@��B�{T�����䛭���`8@H�Vfv��h���^a���Q����S���?���T;�Q���/Wx\O�=�|�e��mc���yGd���G��o�%	�tg�j]�z�)���p1���/����{[�<Z~k:�u���w���������7��S����4����#«�?N�&���g�������CZ��/����T��ʩq�����-��7 (��C�����]��3�UO4{�ĩ-.�2b�ȉ�%��Xڳ5��^���^�������g	��=�cϪ|�Y��ypG!0)�K�����+�x2�w'��=s,�]O�A���Խ���?F�:5A�C�ooxL��h�t9�q��
�������5#�����i�p5��־�.ݯMQ�͂f����_ѭ�J\t@W�~�ϵk�O&��jq7���]��u}J�S���0z%<hJ�i\e��̏����?VS����}�aIVE�0�)�\�z����}K�
�nZ����<>',�%:*�Y�\�JB���*ǚ
"�:��E>��Ǚ�	B������ʁ{N�0:�j�/SE�vf\��'�
�6�w�s������ш��y7MO��zV�`����_��PQ�i0��Y�e�>̗%{��9�
�S�,�nx�9v1	�?sa�/�-?Z����������}zI�a4����B!��4X-9�ل�熠�%ɨ��N�׼}���Wa�Bs�	�5v���߾����(����'~�R�ݞ��'�]L+*�}m�b3~�]c/�o�� Q�.$_X,E�怳b�,�v�ڄ�*���w;L4�R@�R\�[�;W���5X�P�n�	d�A�#.:���@�H�j9�f0�U
Ii��0N�DpEYN*Vć�{��HV��S�\������J��%AҚZ*B$����i7_���7h2�� �j�	���_W#$1R�p��7o�;<�&<���/eN~F��V� ���xg|
UܼL4� �Q������	����="s�w{�m@gO���n�:���_��Ce��C\3V�d�m8H���@ĶO?�M���d�[����ze(��A����r�O��<�dՌ1����:�����*Ӌ�0�g�bR��e��%�h�#�ى��es�|F�����|�_��sU	�!�?J�z|��t�@�3��cZ�e���:C.7u��ş���΃�A�� ����0�5�
QHS��) �X�I`��Z�2���)�ggݙ�nWk(`���>�0̷�Y��}�-T����EY.InO�k'f��!��~=��������o_���m �;kz��'b7M���{�'�#�ot����D2��E��#��j��٩_�Z�XM�h\��D�u_�rnu�"�4g�!�7�|qY�
�Y%8���ｺ>�F0*J҃����v�$��%<�fW.�'�/ú�yl�XD9�����O��6.)��(/ݗ*���]�s/{��r��,_FI�#�^aYg�������r`I�R�	!5O�`e_	(��ĥ73�}�]��V�~bNK��q��EIW5��_ϗL|���/��}q��+ L��rхg�.Z[���-��/�lD�VsZ����*!-�:*���. _)X%ɳ"L�(�'N}N-xp4��h�B�j�)4נ�����I�Y�碭� �]Q���QU$u�B�=[�W��'6�>����̭�9�{�B	s-�稚�-��e�M��c��Z��N�[}_�[�<a΀i0����6�l� ��ꃆ@u�n`^�A��g�4_5҈�w�&~I���hsӏ�>��)����,��O����PZBc�O�w��xQ��{ A��$ձc�'��tݵ{D��0yͪ}7�i�\�/,҆'������8PΣ�i�x���pM^�Q��8k��qi�sj̡.�Z�nS���4�*�J{�ޥ!/?���Y����ӟ��zܦz^��kT`~OO����j�N���1����-&��*zw�{�8�z���a.�[�uQ�d����`e�vت4�H|����i��\�)�,�B��[ 5��A��r�-o-"�	��A�<q �:�L�LL��ڊm�e��Sf���朁%�o�*N����R"&��B.-�ӳ� �	�J&{�����@��p6oj��W�R�yx��	����Ul�g�
�^p/�|��bȅC	�x�Sڬ�J��;�a�.�CO�����vH���G����o�����Z6>YW$7.�>,혇�j�O���A)��9Y���M�f��|AP�;.$���.�n���bgqh�l��9����̹�6�k�b�j�`��mNc�p�Ϙ�F�*ul'���N�[)�,|#�d���K�NR��c��r�йd׍�V��	���2s��Lk�j
o���d�B7�q��T	�á�1P��4���_Tt�&�L\`�o��ox��UڶxF��/'�k�g����챘�bR\��k�zB��`�`Ї[Ok��T��r����H�H��(n�O-�h��6T��a�����P`�V�n��0.�<+�	/���!��Rw�pW��j���Ƴ�O9��;�Rvr�3��QQ'"u��z����3!	3�k@�8Dw�kcf$q����o�	1��N����R��W�O�7[�T�,���Ǻ�lV�pF�j
è�yK���aQ�T7��X��*Ua3a�<+)
�=�I o�[���z�*}� Wr.�r>l�w������"�QQ����޴Lz�6�H�)�\\�s"�U�(!r��5��	��x�S���w��aS��ӓC1ܚT.�FjI��}��²cg�5��=%�,�C��?"�El7ovJ�v8{3"4j��O[�fj ����~;��=�͘�-K\�#%M��;lDN��I#`�=�����w7�j���1�%`H��lpZ����]z)�*r��!o4e� 	��4�$&�c8e8����0�\�S	h�Ow�L��V��/�/�\CUI�
A�����ZC<����<l��w5��@�"��,�
�<pQ^�l(tH�^e�q�Xs%��G�<�ma��U6�hE7�7����A���C�u�-ĸ�r���:��>+;��F���&�	ïcQ���Z��;藡��/�Yx�e��9(��,� ��;Ea�7��X��~�_���n�wtN��(;Hn���5#�B|
�a�^���Y���OP����,XlxVHYEB    fa00     700�k� (�-6��*E���p��t�����w'.�M��4Z�0���[u���m���`/{o%���:�>F,"�+�팃M	qw�|N;��� GD��7�O��H���5����I�@�)H;0��U�Ws9Djc8�t#Ͼ,��'a�k�d�)].�ŵ������Z�z��!�"m�wB!o}���oT��u tG�"1X쓪]�� ��L�r5A�d,v/�)��{yI�
�"Yr� uy�8��1�tԥ���z|ot>�0�q�J�#���ò�	O |�w,�O�~�2������/w7%x��l*�K�'^`��f�����ѽ�I�S/Jd����Ñ���� ��IbyPTO��,�mM�"�kl�M� �9j��H��j��G��:NVw�Y����KM�����d��;nw2��v��0��i�Ҩ���ؤ� �����܌��ڕ��88� ���W�[زc|h!8Y��u�zʸ�!J�0H�e93��9²�/��d�����I�#��� F�C���m)�Ŋ9�r��0��,ED�V��M�T%�ΛSGw�m�'�?�jn��"�mX%��C���(<��L0LG����،�G@ˢr�=9� ~ͪ5/������QTr6^)�K�Y#��qϺ!���� 8�,�n��
�X�<9����i}���G���+rЇ��Tp����}vD!���;��|��ov�V�m��m�D0I���z5��a�71���#~�uf��Z&���LE��K���|�,��f+��4�^�&���L��-I�B��VJ�jN.�|���e�?�h��m*0F1oC��k�����z�H�J֭LEe�:����&�s�`1}ԥ٨W6�Zw�*ؤ;��{uT0��W%c�����mi|{9"+_	s���ܑ�A�b���#.yզg99��t���֙e3$X����^}�Kb��w��q�ļ�w���"͕Q���/m�ф�\�P����]9�n��AN�[�0�T�cL��Y	L�a3C��8��;8���A^�͊PC�]٥�˴��M���Lg�Ѥa���S�&��q �[��}�½C`��jCD�	�5����\v��kBȧR�XQBz��w��8����x<^W�������'L"8mZ﴾��'�X*�H}�.|ɠ�g��5r"E���#{����%]~�
�Wa�w��(���B��7�wNu���Lx%��Ōf?T�L�PN4�̡A��&�<�΃�&[_��Kxl��f\�h�
�33���OG��0��(8�:�?3��Y �0Ib�!}\۴nQm��7M4� �� �_�-&Y4^b����*6L�-����ub��*V�+x�t�BCIL}�c�"2s�(!$e:�1�6�z���i�2��U�.��+p��ʚ/H#\���2Ԥ������>6�L��h̽��;�;��d�EZl���$d�~F/Q���TrܴKE��V�a;" �(����sӷ2����=q��}<{~�Ƿ���lٔ����ݡ���~��u�^_�t�����:�l��q�*�Ik:���n#�:�d}yUU�?8�#�~|0���{u��+#�\E�xp�C5���m�̺a�P�I�.`�'��Y��V{+1�ucą^�l�I���z*5MJPaUZ@=Q7���]2�9��0/85�x[Zd$��PȊ@�#���/"y3������.��	p�����b��4+?��%��֊��|:���8����Q�$=�!��^�}�Dl[rg�J�3O�~HⅮ����i��c�G��XlxVHYEB    77da     a607�a�f_��AV^�|�G�(7M���Ub�xU�h�@]K� Z��I�j0|��ae$�1Jm>Y�P���M��o�]���kw�,����6���WN�c������*7괝�$�7?;�r�ɢQ����͒�&p ByF
�xN��K^�1�J���������>U�	~F� \q��������_�I�>0Z����'�s]���Q�vQ��7�Q+.ng�z�Y�C�,S�yyj�$��c̷Eߚ}!���G�qT�OB�Mɋ\a5���f'ψ�z����f����y��>�gr���%
3��R��Wq�L��)#����v��w)^{2���?6������.��b�j��F�?��]�-�G�h�t�b<�L�J�}i-D��CO[M�{J*ޖ��ć�`Y�8tOvpN���0�meR�l��!����B�wTD�ꞛ��c\����H�G�]z�̈́z��h@%�A$E[N`���Dy�H��l�WE����t.��P��\�8��@lʘ��(�Ai�@���\�����$�T>C��ᩕ9��Bj�ZW���n��	�/ߵ�p4�*�8���������J�Cl߻�QW�
���ז��j�8$��m���z�k��GG$�����?����U3�Q3�w2]�f���pa�;DY�{_�β�S�:�ZA�����kV��.�{-P��PwsI6kֆ�����pZ� \�UJ�"w�?�Z���!���X����I�+�e�Y&��A��c���lN�1a�mj�3(�zt~Q����ߤ�\�T��^OL����6�?���%2�� d<�
S��­���;�kۅ.�z�����{���27n������
R=�*�٢��c�c�f�ܴb�#-���6�O�	�<Fs�;q�S`��]��	�+�&�
�Arȩ��gfI*v+)���z\�x�ĵݵ����}nZGU���J���J�#�_	ɟ�P�!';�P\���b�˰@�

���־!��5�;w4�?	�T0l��B3�C�N~�������K�MC����*�y�j���6�MHe�E�1����� �R�f	Z�{�	 \	�C����Z��(��|'����"�%M�H�Z1\�����a�A|:�:Z4��n�@!��J���uK8������C�\���0�4��q�\G�����1����&[���Ք�-8^���|�l��o�Y�.W����z��I
D�a�5�.������*�؋w��T/�H���G_���j��-�e�\�0m=ܿ�E��KJJ�}����H��3 ��~iY�����o`�d��0c��k��%?�C�jA��L�d����/ x�!N/�v2�)׉�M�|��{������>���ޢ1��b��[������S������^e�fM�����6��>JrJ�����Xd��Q�4�4��o�&�|�'��9*N�e� \9g�x�j��h�?� �+#�e�K�Gx_c�e4ʚ8Q6LtM�*�o�D�N%}�tUeW��ϯ�MV3W��[��	-;-�8O�Н��:>�����T;}7�C�U=f�A�b^�Qb>!���B��2c�g▹��?}3a�W1���������t��y��LY�P8 +�߈,�)M�Ht�_���|��G��]"y�;RR����Z����	J�9qe�3N� rV^�>������)f���T0�5�}`��j�< �q�AO��L3t�� 0�� ��8�	b�Ճ�f�^�a����EW�W/�'O�@��e0�EW�?�2]�S>�~�[�\(a�Hԝ4Z8��]�X��?𾖬lfw� �\5?����\I�P�Q�b��s�Z8��L�c�/�1N8�=�ꧫ*`rj Y�[���eJ��q�[7�A��0Y�D<�z�Rk����w�
�H���h9��f����b2)e��,�F� �P�N��95���ǜ�a��h�6:��Kt䩿��3��m����O�-�5`R�$`k�컑{�C�j���(�@�@,6��].⧅�,D������T�V���2l��Ҵ*G��L�Ӣ�/%�go ��y�<���B�4�1�K��fA���8>,��i�t0�Ͷ�~�e��d(19�+��¢|����%����$E�=a#ɭ��j�����őP�<3Llؠ%�����%�I�̑���t�n/-�w09��R������!Z���Z�����	�콌��ଲc��V bf_��>=�b>��~��x?�?���o2�-��*���^_W�6l�rֱ��v�OY(8�sE'�w�K#ߍ��,�9��里nWSĚ�]-a�h�I +���	 A��)����d�@/���Luܷzq�*yե��>�-1 !`�$O&a����8�?�SF����#����gV�����ӊ�%X�GM"��y��l�"b�w��;�X�x�ZT�*g��j6�R�6�/��y�b]���ŷL�,�[�9�<�]OAK�h���Qb1.���@��/�o�7����]<}YDt�ܽY����M���ػu9r9\G����]���f���Hg[Sxf妮�I@k��k�/PN������l��\x���;�	��K��x�������