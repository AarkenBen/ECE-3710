XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����u,@��M'�=/����ţ&�-9�1Z��H��IR��<HED{hp�c0@���b�Sm=/�͹2������IQ���~��W��n��j��w�>��2f;���޷w�|�d�1���纟�]�[_�3�%ᐪ_���E�>��'�إ������:�ﴱϯ��O?k2�sX'��(Ć�፮-�H'���
 |���C::%uiӚ��{���hJɣՅ�~o��7�h8�ZI���Kє�}����;�nG�*����h�L�b�w��D-c�V�����/�a���i�u⹒%;��F�^dԟ�=�����"�!�d}���Gɼ^�j1Zy	���l����F��F"^Lέ�-��8�vԀ�5��Odt�Y�mpb�f�os)L&��#��[�4i���L.U�7��N�����B*K`F����a�Z�w�?�� s*�"K[�ZT��3�����������e���[(�"��i��2�&s�ۄ��� ��,�v
%"��%a&����~=�%Z��F�!l�ʹ��`9��vǇ����g���Қ{����| ���:*�9D�����ھ�yV���X��f{n�����nVQ�8�sa}|�hg�	�j��*����)�5��}� ������G�D�g��m��L��� vKutg�l�{��q5���f�h�g��g�x������٥4�r�]j��ڐ�K���B�uGo�&|��;--!���WL�.E�~�7ݴ_XlxVHYEB    c763    2600I���O�a㦺߷�# �Q"�0��.���U
�$⍽��Y�B�����s���!�J�ܚ7Dy�U�x��*�3~eJm_���aU�>EU�so�>�G��EAcJ�N0�&g]�B���`�Q~=��&zʲ��Q�MS���/��l�����A�PB�}z�-X0_��^�-�Kbx)��Q7��W���y�^��8�X�ESM*�1C�C~tX!V�5�� ��@��|�mr��t60(�o�R�G��#�� ��V�h��jkP]���� ]��M��,M`�L֒)�X8��˺��_'���+���Zl�o��"m
(�5�CyDi��AJ��uF7���VF�CC:�\G���c�/B��bs�����lt�>ie)k�؊���;��	[e���a�<��x'L픜2f�2:՛dk-�]���&2:��J����m�?��Z&f2�I���Z���.��<ό����<���<��6i�7�a�=�%�D���5��m�]�D7� ���SV�J�[#�Hd�Q�mMT)"7��4t��:��8�x�Y���0�Gv�ݿ�CU`}8�U,�p?:������Ƹ�K��J�3�_4* �����g�+@�m���{%�G
�X��8��}�k4�Bq�)�2e�� �w�dv��o���]sg�x2[�_xL��!P�H�B�EDfe���*!����r�ɝt�A���7���݇�J����؈��7c8�!C�j�oR���2��pD�2��J̵;8]�&�s�{��(1�����;;�Q����ߘ[N�axk�Գ+;Z\(�����^K��9׼֫���3x�mϏ��J&��a#�}��ϩ���C�k&�(/��ݩ$*Z���Wğ���j �u+�yH���n�闦0Q� ݺ�~e��;x�C���_������qB$ٞȃm��N!p��  t�'��@M-�����p<f&�� ����4Q�ZX��`��%��Bz-N<]<x���iD�Jw����즒 �\�Ѧbׇ��_�����A��,�6*쁽�����"2�2��*�I/w:�L�i���2/�R9�3��|+D*2_c�vTI��Q ��~�O��:<�Ů�)t��F�����dK>�� 35I��$띝=���`T �E����8n4�YBHJ�P�!��?"A�DT�BT��Dty�Ħ���l�a��9'���jb�j��R.�LR�\���Z����T��/��(��$U�1����!gں����|���]2ͬ�S1��2��͖�u�#O���˖�]-��aV t���*h+T����Mɭ͵���]r%T��І�M�'�z��]5�����~K��D�Q43r����)U�܆�A/JTA�����2���ʾ��=���M�g���>��´Z�Ѹ��c1�;���?�����L4��A4�(��j�w�}�����a.��g�EFv�J+¯��fhaB��L�5�e�&^�1��8��s�k���?���~��rS�o��y�&W3C�0��#�ۂ�9���80�<X�ωP�]�	?M�癫oZ2d�=�,�N�S#=����T�2�bM�f���qf���z�gb;c�ʼ6�ܼUq,���}��M'����P�~�Ѕ����\�1�&�d[��'ϭ���H6���`�gOj��":��<fZ\�vtV��5E.�墂]mS�Iֽ�a�����g�]��.b����6"����7A(.���h�%�!f5�(�q���kM�횖���A��� .���TG�Q}ÉO���{2�\�}2pR��]�G����X��w|c�
t�z�{����?.R��ـ�3$6�V�؄]ٯN��M!c"BeA��d�D@(*�3kh�ymG��R�����2L] |�3Fk�g���[�q�v�����
t��b U����<~Cyt�I��k�^�V=k���E�{N?��ӈ���A/Ƚ��2XRY2T8�O)�үӏ�y=K�)Z��a�/j�޲�T�OF�&×��쉽��f��E���S�C�)��W[**�j#�?MM7�G�v��S ���� k8�I8X��uƂ��Y��T��C8Jv�=N��h�j ��ID��쪿��@�kO���1�`Gc�q,�Os�D ���0����z���I��z6����@sf��Dڎ��<��ƀ�rs4&�5���
�h��(�l�m������vO�^�/!� �*V3�yp�NrQ�I��Raz�ɐӕ�,�\� �%��$�s��C��T�=	Ji����������Ӗ�%;X�;�\��^^EQQ'	<$ev�9)��9�g��xl�vǍaH� ���u`M-�S�B��Q6}�(���My����=󟵑�ޱ�S�O�|%��\��)#�=�`/e�'� ������:��U�G��2O���)J^ԃ���=\g�r.b��!�_�s�U?�	lF���K%0��-��
*������a���SÓa�cR��Vm����f�mi_snS)�7עLz��n�u'�u$m�������A74l)�:-�Uk��"V����@���RIm����F��|��_sIGg\t<�3�\kt@�7l��Փ����ق�hk�f���q�y�5`��K\4_���H�����a�lD$��.ڛR~�'Q�&��M �X��oh"�v]b��䀆��(�B�/�!��m^"UxnA�)@�yO������E��R`V\Oo(��<"�Q-AM��}�;
Y��*rD*М"�y�~z�	�ZR�3W�)p�_�g=-�Y\�,ё����*VX?$�'1�=�v��%h1"MT%Z7!N%D�Āl:�2�a7�_2�Xb�����]��Jя0Ozň��;P��e�ߴq��*X���oP�<��:���}�)����!:n���u2�0oM� ��^+tV��ҫD�YRni���$��&-'xA������U4���{<��+��k�fӱaqY��Q�4��F�'V��ն��� �<�+*}1 ��Z��Y?��!\%~U����W�vC�z<���ܳ���;��=��,$2�1���Hv�o�ΐJd�W�D	H؍b��/RV.[	��i	�8h���m&6bL�<YJB��C?_���2O���\GU_j���VV�5��8b39�j��="�(W��kv�":�~結xj�[z���q����j�Uk�c8��i_�$�:��ֽ�$x.Lu<�MYg|���}����ڬ,J�
L��k�a3�i>��4��NveQ1c�$<H�ύ������6�}�W\:�(+��������'��'�olWG�Tj !�a]�$'�b�E�5�bن,
�(���T�zy��UQ�!mc����U�bQ$�]֙�[QuN�7��5p����@��d /v��`�C#���"��c�H��ٰ"ф\��VU�6Sҫ)�����oJ�a�}����~/�<����rF2D�:I"d(��#����^�� i�_����A4o�}x�O�"L+�H@s��R��2� 6t�rP^V4}���,����Ȍ��_��\d,]�J)��r�}X�d)-R����L
��0;�}��-��1�m(��ï��B�j�����K�c���F��X�Wy���?�S��2Q&l�N�(+����'���/�{����$���|z��S�\/�����b}9b����ySW']HY;���&�a ђ������8��c���)�8�ss�=��M�Ϡgo�MA��}`�8o4U��PՁ$v.���Bz�L��Qs���衳r���S���mi��I3�)J�Q��2�~nϬ'ڠu���VW�O�úCRu�	��猆'C��	"��<6+��f�%�]��x�d.O�%l�n|e�[��$��$}��ߩY��3�¬�J*7�ǫ%��%V~�Z�<�NN�b��o@�l��:OM����G�OTV<�-�=F����M]1po��*�蓦�� ��%#�<���_;�~�Tzk�,i�h�8��:lV�B\J��:�}���u�D��x�u�^	G��1o�<�F������ہL[[�s�7(��i��2���g#�ޛ�U��FZ:	��͟b�YH�.;��4���4 �����$��ƻ��$G!G2]�A�a��.�t�5�� 8�Ȗ-��<���/�����y�m5O�𞚲��E]?��8Π�L߬���s���0I� ���D0���Q��m���+H��Z����Tm��{�ٕИ�v��(����u֕�6����Y.C�N,�3܍�15\�dXKCg�J�N��L�ď%�d�0=&��ϣ�z�Л�/���vr�.R쨘��{��C�c!Dӣfq��T+�Nr�]^djv��01�z�  �GTԢ��=�
������;�k��A��͵�b�K2F�d�{ԋl�T�p���P�S�*{,�3�ڤ%>@�9��;+.Y�^�ߎ��_�U�����K��t|��oݜ��]$fZ�ytf��3ڇnH����LU��I8��F�$�Fc�-�W��̀[
�F��bM����KI�K�W��7=���</.x�9�;i�Eh�\]��4c�c?ΩN�$<PG����JC�}�㙨�l��8r��1��m-�y�!G�������;.<}���Y�(��S�;tr�jw�M;IJ���7CYG��-ߨA/z��W�y�s�X��b�`��w��m��\�zck�B���N:�x��+��᳥iJ����)��e�i�Z5��q(�R�w�y�^�E�aAR��71T�Q�� Z��w�Slܵ>��v�FPh?�X��(����-�d[+Ѵ8K ���g� M0
y^�U��Ca;1!u��?2�iӫ���y���2��,�}>A��>���MS|=�Q��
63�������6k��L�?A��4�5|x������.ߑ��v�¹�0�I6�,�P�d!��W~y�4�G�r
�7���ϺLj��Q%���}�Ӱ�bq8u��3v2$����5� ?j��.�~_�����k�����H!ۖ�>���P��s$/����Z�E�g�����Z���G��fk �:l�o�)��Z>9���� ��6X���?B����`�������&>�I��#�`��I�>�+�!1��ؠ#�^�ҷ�'�I/�.���JT�^��=Z%c���D1�q$�Rv�����1(�3"R!���E�"�i~lW��z�+���.���,hy3,��md�GJ�bO �[@�/m0~	��0�ڵ�����%�k��`�^ ?9�c����>��9(|�_뗽�'lq���g�t����e�������F��.��L	 �}�	4D�c���o��f� 5ԥ2�ñ��\�Ck�� ǂ�ɐ�J<}-��Coy�Ջᙼ����%����a5ȧ+�5?�.U����Z���-U��I�&�{y]{��h.��� ���%���o�PB�!��л��e��^�|�R��RDtl~����(���R��DG�{��R��xR��v�T����S,���X?"��ȟ�����i���2�i4(�T
���@%��7��	�*wE��x��6Z5g��no⬨�[��a�b	���&t�~��e�%�Ppu��pC�2߆��RJ
�7���K�vd�o�|��0b��|��~�B������eu%u\ϑ�o��;�WYv�w�g1��7��h?�I͵�/���G�!5&�8G��z�0_1aV���| �٭��9'&��k�o٣�A����.V���.F���_W�I����O����J@�����Noō�Ph��C�	l�(�;�Ħ�c5��2i��e�`�c�g큕[rʍ/��Dӳ�
d2�+w6�����E	���o��]g��LV�-\��.��aqڤm�F���n�$x���a��mZ�G|��It#��Ѽ"��wD���>��v��G� �6t�cݭ���J�1���'%9k^���ì�k�g �1:�a����e2�ӵ�f�)�f�f܇`���(�cU)��M
SE"r^zgWu=��+"�|�^� ��iL���4IO���h�"��A<��5Q_ٯ�\�%���S��oN$o��m,��`�O� �[�1�3K\��&�5(O⽤^�ʪ��.J:�9ܪZ'���Da�-����A�hH_~��>�c���bu]�WEPD�3Ӳ@|� ��iW:��F����U����]l��5s ���|}b�H8�S:I��(�f��i��ʵ�*��(���n&U	�_�*����᧦9������ 3f�l�g]dv�P�qHn�Jܕ;�m��qQfb/���i��~)F5�����RQ$x@nS��$��
nky�[x=��)���/�����ṙ[ܞ�s������A���š�hA8 \��욵P{T�Dx��}O�d�p���S	���˲AOr?��z��lX�'���!V�j/�d�>��;C.�_?�������X�!0�8<���S������f��y�R�m��(��?[�W@�V�F������U�j��Zo��F�p���ÏN�������*�����9�΅R�X�f�FQA�i
���J�<V�)��������	ʊJ����Ǣ&U;&#�@RH̩۲���9� ���� ̙0��S4�ž�0��p��5ڸ �2V�>����ef�}vu^��%�r�����\��}���c1�=�&X�Ń;z<�j��l�:�~�{��K�U�!�����D!@j`J���U��3�Ă�Wh��E/P�Q�-���l7�n�ʀ _>h]��n����E>�*F�����SU��C[�*�C8�7��e�z~�	����7����I����!��n�l_�#,�d�=���$�vb 8%-�D�*o]6^ ��{��G�}�"�u}�w�s~�؄�6�3��a[���#���ոs=���'"�=p?�:q�?#G��6_�qX|��_jZ��e-q!��@Yy``G,��%+��;6�hU'%��G��d<��0�M`�%�x��]�MqqV�����·iZ�Z�&n�P�u���e1���ǵ�i��̯Lk���|�/���	Y�n��ܼ�v�ޟ���������?��-���W�M#��A{�w��6p�M��Ce}>�e 2;4i#q�po2>%f5LA�J��9����9���>q�@�h�X�0Z�R��f)k	ϽL5+L�������v��TBD08�z��U�s�a��I���p5��>�s�kɢ=y�i���Y�!E"�;%��A�V!��#%A���!v��_u�s�[�ꁯɯmfXd��Fb�-�p=�c=e� 	uIDj�=ͳ?zmKjA�}���̫Sey�(�h�M��>�B�8��l����l���s���s�Dy����~ޮ��G��`�޹g�aų) �O����I� )�){R!�)�� P^yt�B��g��w]n7��yA��!�[9�C8�V9t��㧷��긇Z����b{�J���	���o瓳�����Źk/xs�����:��n3o��G2��V#A1���~���_�?�EU��;����ҝ����.��N*����=������=��d�x�.�p\�};���f���l��$,�2��x��@��׿"��4��۲?_]j�T>�D5�D�b��NeDD+��y	�;�#�^����N?��"�Ձ1��Ot�'*��jR�y_T�6��CQFX"pP��%�I�Y�p����F_ԥ�`Ԁ�6.���e�a��7�>��n�;Ō�T�Q��`���m�B���`l��J6�:�B.3�"��;�A�~-Z�y�G	�.+p��]�&�8u�S=H��O��	�*�T�-PSyzK�NpM��/�뱔���O��$������]�+�	���j�]Y�M��v�ި62���\h����M�?���#'JN(�5"�]�]�
r�=��� s��3��&�M�8��- h�d��ێ,�.`B㝨��\}�Eڈ3�(M͔0�H�f��ā>�m!7�&�0H�PN�
8"P�҉�+ٔ�W5����n����+�) �W��'e�"� ��D����EF���n�
���Q�6��D}��X��E,���f�@���͘;A舨W���Qfj��v����0V{��֟M�_֫��ìo/p��Y3j��Lfpm$뙽����wC_�|�k��W{��~@�@jcѻ$�41X��p&��Y~K�_U02<��ǅ%���Xal��
�q���xf>K�|��[���pJ���%�r���
&�#��BY~��Eh�f��Z��{��w�����I|󔳠�V8�ff�{|��Q���o���쌘M|Y��GD�n}��"=<78�!ҽΏ<[$��0���ȥ6R�����(eU���-y�(�8��-`����wǦ����)��`.�\ZT�\��0�3mU���T!��W&XV����Lb��&���[Dz�Ò&�Awf�	�>$�n+������o�K;���H0�K�B �(�ƃ,�Z~� ������)eT-�XQ�ˠ�9n����_`=~YL�\k�)�_o1��O�*!}�N�H�>��vwtw}ud����eז69"����:����rr#�l�&���&�#�e����<��q���k��Q��S_�>�E�Δ$�D��}��cT�-<��$�s�#�����wΎ�ɂ[�K`1�ڪiJȶ���O�Y���7O�X�����a�/�e�Ղ,�i;�[���(�Z���lH���G�f�\=Y�n�w�-��ZX/�'�7�}B����p��6p����mp���8�ۂ�>*�O6�sa��#ƠV��NQ#����P�M����]\b}�%��0"�䫤ٙ��Q��O%���]��ز?�����|������N�ث�縹��@S�D^���y���1��V���&4P
�-/Q���{6P	�X�T22�?�J�wO��G��H��sIc!} *�]��8�.��$|V��HY����ŇX�������̣���S�.���]�DP�*y�eo@�x�rȞ�� �q�m� ��Ȥ�ZaR��B�Q�
���PJ_���Ck�'����D��.�Q.(,�{?ſ������(��Km$nC��̞jeg�"�J���`���!ޜl�oL��ݽ	��y�����z���s�(��
x����H`��r�n�� �xޗ��D�)�g!��O�Xg�1�Z��T��}m4Qc��Zc/s��QB��5�R��,�O�rs�K��'|ZK�	{1��|yq1]�zC� d�c��R�
���`��'��T�4�l�j�lU\�n!�@.%����;��؆m��0g�,7pqv��l��=z��X��[mCR�-�+jb��Ҵ%c��I)��x��8e�g�&=��@����(ZS�f�dT���Z<���d�6>��9p��d�P�o���ֹK���*�Nq�cw��)�CI
+�ۥ�{��^ �����}�hZ��Nv�)҂��Q�TNl��{�9/�����&�5�k�4�C����m���i��O�	H@������Դ�v�t����n)�`����{F�i��2N�