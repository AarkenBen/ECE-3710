XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a��s��Mײ����D�*AŲm��\��Gy��U����;���Ϳ�������S�6%"}����Y���eLƸf����v0�����i~�eA�\"v����_�����ɚq�c!_���>��\O߶8<�<e�����6��Bw�?����i��.6����ҫ'�t���ǡ~R9ǚA|��������P��h38L���pHD1�uez�� r�2
�!�(Ⱥ��7�xnPGv�WJY���~b�!�rz�d
b���y��zX���J(�9��|[NIÈ�����j�;x�/�F�G"F:0���i TR<�~��Y��Q�����$t��*�W�� #�S����1tC�B�+��w���/�D6�������e������D'��,���M$f^?R`�;gk�7J�>��V���l�~��]����nR�
%�))�rj�Ȑ���O9]��9h����>��W)i�q��״�l"5�x�^-���HIb�������� (Z���c�qr��+�D�g��0��@���O��޾}���#�Kr�I,��@�bb��G9\'�z��Cy��+�'���.��S�K�g(��L-�@c�=��%��	j��č�q��{Ń/�ysWCDwɽ�:J�&H����]����I��h%c�ɕ;�ˮ��r|�6��0x�R�~��EX#s��n4�D�6Q��M��y�B��P��+g,*�g�b��7�}�QB������A��m\�b�=�)�XlxVHYEB    29da     af0t1���q�+�=vbf�VZ����!] ˶��#`�f�=G����%�f~Ԋ�� `qi<a�NI>Nc�D@ή�U�1�,�w4�093?�&F�ò�?<�h�@��]�$�9�gq����r��ÚJ�(]q�K�bU����`����LQ�V��C�1������眆�F-<��ݙ�'��m �����r����W�D��:oqe�������b	��\s��o�-K���K��@�d#>�fR�� H���z|lO�,`�v�ֶ��9�X��-�a&�/�gԃg�Q*:��zy R�_�]����zĤ�C�cӛ�l��v,Qi���E�*ۏh�ӠZ���.PǙ�m��d�'�����=�2OnK��+"X.�9���	��:�Ժ��e�ʦ�J�]/�!�1���ZK蕈�ۀG���*/��h�}e�`�aZ�Jz��L����v7����^��d�IMR!��MW�6ؐx$.RUL_�c�QSP�I|�����F��-fI[θ��$Yk_�XcKzJ��3��e6�V��~�*ƣ��6�RaQܨJlĚ�ߑ�T[�G2��A������}�]/�iuv8g�!L����u4����Ǩ3W�Sɜ ���8u���N[���0����<NL��Eo/RX%8��hU�/�{{rk��M�ܚ{ڨ�C���x"ژ�Y��#`Pz��"R@]��\��n8���s� �o&�%ݟ��6ׇI6Xx���:��;�HMX�:1K�]XN�C�'��`�n�"�ҷ� �)�peʩ��=_��r�$����M����,_���f��VK!�:��'b�yj5�9�	�君0�L+����L���9��� #���7�Q�a�ܛ��R���2?��~� ��U����Т��(�N�$�b�"� �P�M;����.ή�G��_#.����hn��Rubp��I$��p�m�Ic�thǎ�?,��RT����aXjs��?Q��\t#�tRn��弛h"���<5tT�\�PΨΑ��l���q|_�n��+Z�,��Ro��C���ߖ�wj�"�8K��@�C+�t�"Y�aq����K'a���zб��kYu��L�-����|�
R��p�Mt�7*���b��IxX�h�/��V5�d���х�Z�ޙ���l�P��&4�hgw�)t�Y�(��7��׈Sx�c��F����Y�Ƅc�	:� 04��q�c*p.1��t~0Q�FK�+.��CW�\�0�K����p�� ��PO�x?0��h0�?0�pE�m�{2l�g|�O�W����J3z�鄟x��������p��ݣ7��bt��_�Č�
2�|J�;UhLw�6=db.��%f��R�y�]�aվ��p4|2Z�DX�S��ͦ��8���>��LGE��m��z��X,���.1&Ap��B[]�lo͍�WA�MF�L��9��fw`�� ����ClPSY��~A �t@�G�<���>�._��&�W#(�k��ym�
&P�Rm+���I�di��#�@� ��Z�*O�WC�1>)�m���OnM(톑g��DY��h[Z�x�qa%�:��cN���e��+n{��ӧѝ��:�׊"�hG��;���e��R=��Z��~,�[�n� �Tf�����݄�I0��@�6�����a���vY��v�����s���� �q�[�1�Z�w��;嗩m ���ZB�H�H�V��.�+i@ �+����(;��b��Y��)�e�}c���	[sS�
+�J�U߈�be�X�ꩄ�U(��e��	��FKo�q`��W�I���L�,�to��W���3�W�6!�G|�)i�g�U�1.����W�`�"˥��2��D����{�i���'�G�a[j�<1S����iѼ��2M��v��+��&D$��Z��E8xZv-�Չ���p	�����`�	m^�3ry�_�\_�C Q�4/��g�П�I5��C#QS����'`��k����xW���.��$��M�m��9��fL��������m���Bu�uڥ1@��v�o�'cD��
gw1r�8Ǐ��4=��������k���vO�&�4x%�}���s9�yZ��.���M�z+oG�ݱ���-�B4)i6�0~��O�C(� �ik��ʗ T����i�"������__�`M���m�k��N�X+C�=����)%i��14g�j�,�R�m��դ�>�x�����!� �(n힠v�]ڊr5�?�?1H�-�Z�1��\��)��1��6(�0=���x��4������ ʋD,À�mYw�ֻ�d�`�Y?�㗢�����:6��<�N#��Y�)��2pH%��^�g.2�����Ȓp�O��!4r8hb�3w�ht��l�<�:�>���_S���0 WE����w9�S-k���{��RtvءN��;P�`z��@�c�ݭ/���h�$���{ԋ�ۣd�8NO1t�@Zh���=�x��.�R�s ,���J��������gG��s��"h��.��X�|��<�<�+Q!W��'5'2�+����q��x��(��ק��ܒ%#��h��t�pb���E�u~@5��O/M�o�g,�,�n|-�!���#��Վ��a�M��7$���ɭ�A�v�w*��	f� m�8�]�F.7��%�)\�o�^|�-Ot�\'�*��^��К�C$�l���p���By�y�g�S��.�|�����g����3��>d}w���