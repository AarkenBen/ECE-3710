XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T I%1㙘�;���-�'����;��=��s��._�)�͐CI�`7 ���E�|�{Ot�u��&Ak-�5��.uv���z����[NΊ[��/a��1�=�:��CZ���쓱����7`8��_g��"�}��� =d�������M�j�u��(|�������nQ@��|�⠠��FJ� W
|%=�!x&Z!�~�mhf���-�?Y�d���o���d>��_�mO�e
Yy���?�>�kqZ�/��{d�%ىSg���!Z���͗jf���W��,/��x0u{Wz7���V��$���J��
|@9H266̂�΍9��W#���|X�����)�j��7K�)�k=ah���^4��|u[�N����s��p��BB�K-�g`��{w�,���e�[�G m�9���~M[�)�>G���W��nVF���$A��f_���,ፐ�m��k�{�Oenu�l�q_UV�[�$��L���� >�����Nlۏ�����e<�)�]��$��d+�ؘ�5���券UD����
��fM���c�UdK6E�Ǔ�{��KY; �(��8j+Eiɭ=�A�]k+��ЧQ ��"�e��W�[ð�������#� ��O��S��l���"��fʖ�G�V����"��` ��nQ��z������B�u�L����QE[Fm���#�yUԡzgQ9�v���	�:6fk矴/!�����
�@u넅���Y���}���R�6�-�w3��MhXlxVHYEB    9efe    1be0� pc�t�&�X��&�^V�΅Y�S%���,�T�I�'=�t��*���c�ds�WoN�+o?3n �߲�kTQ�� ���*͛]>\R�~��G�2���vievy��ʲ��0ܔu'��xH�>M�u'�ה�	br)�Q���D=�t�W����6+�IF
(���F���&�oQѬ�TX���s�] Hz'�m{���{�CZ�f{������9@
>�!�b�wg?U(����='P M��t�}w�4����_c���S:^
�/|�B:2�x8�G�?s,���J�^,˛2�cC�������2�JBT&USH�{��S�>$r*�3d�K�U�y�w��c�ȮPEYb苶kG&��e�,�4�e�ŝT������XPg* s%G�Ͳ�%c�}y9�����Ȍv7?͚�| �}�m/)_!�S��l������l��AZ�1��C�rͣmZc�0�|�V4��dj�Ds����ʽ̠��)X1��]�5у�0�)_�D-���N�T.����:�&�#��<R�d�󋗀�1!���_�uC"4!�Vܭ�S5��E�� ���We��)�k[Oo��|9�è����r�����	f�R_�\nt�Z�ic��%������L�-�~L1|�|�>q�L��Pf�`�)�Ot�tsd��þ5��JM����:�vM-5�j�LH#3n���fZL����t�.�G����"�
��6����P��{::&0awql�B	^O�ɐ�[���ŸBg�C���$��}��'�B�dy�y��d;����<��g��8�BO����˷�Z�_�G��<�1Зr@st�/�x[�Vڭ��������{�F�N���w�C���|=�S6�q�(���\�q�¨��s��H�e�>�m���kI0����߾�`�&�1��]C��k���L�İ��zBW7#�����u:�~� �s������f�*�M���W�S��/�.��Z��?u'��z����������ءHxۆ7�n���i+S6­l���� C������]�A��W3�X��_��� �J,��<+��F�	�]��0"vH?O:��b�$�9z�3;I��X%�D���a��Rh�)Y<^x�s��з�Y��kF����fL���l����	z��)N��F'`0k#'
�m�w�1ѱ1����t�*�b�Uu��* }�d���A	K�RaӀ�V�Vٺ�;�[��^�U�ű\v���tQ�L�¹~��9������0���@A�Cnnn^�j���|�� �
�"_شۄ=�ٿg�"d}�2�G�Xc�c���0� ��l�A���0H��4o�� v������ј��)	UĜ�,'�&�j��^�J��=����
�G��b�����i$\�L˓Mg���W���^<�.�7L\�#�JQ�B#Üi��]��4�ݏƍ5k��)V�>���xIGx¡V�y13}��wr�V-n2�
	�O�8B8L�4Ng*�doa��)�j�}����iA�M��7�߾���q�,l5uЏ˦�6Y���ƅ	&�k�)ͅ�wn2ˉT@�H��6��C��_�=�~i*�I�����k�C�dS�s���X0��oDi���l�����w?��mMR��y��
�F�1H�A����mQ�7��ܚT,R�ϳ����ЕCpJ�S�1�?�Kƺ�5����<q:1	p!���#� �i1/�i*d�,�f�s~�R��<��o���ߴy�x������S�̌0SP^�!�0�1��I��[Z���w�N�˯�
lM�T}��4�g�ӕB���I�+������4߆(J0Á@�
c��8��B�����[��p�����yyjo��K����{W��щz���t��C �ñ C�ǈ\�2q��5 4ounUf'��s$q���K 
lCI�ܛd��M�/���6�ڄ��t�p2V�b��˘� ���p	)��ʒhEJ�d5���g+��Ry4#���CI�i��̄�>��|�<�7J�آ�� T�Rr}�ѵm�b�F��*M���-?�Ád��G��~�A���(�ʛ&~���Y��$S�q���¶��H���������fJO�	�S��jK�)A��n� &�K��C�x�e
�i�����
��q�q��r�`��_�m�ݑ�v�B���x�'���<����@R�AG�Dsu����c4e �I�5A(�Yt����6w�̐�
A#9��5����_{y���8�1w�oŻ9�#��Y)���Ⱦ�s�����ۊ��@_q�[1}.( BR+/��4���0,;�����R���UN�(G���v
{����}L��|OI�##�ӫҗJ��'�	�K�mgv-%k�ť{`PB�Zwk�f,�3�ǄN�����Q5=T�����&+r�_4�rOS�����'#{z�K�~���r��fm�Ƌ�G�4r6�D�,TAua+jp�7�)V���/O��SCO;5�T���������J��7����'����E�m	�8��7������
���W`�8\�͂o��)�Wz���
ɼ�	��T�w��V�6%��=@!m�o�%?E8l�F<^���N*F�{>K�!˕a��PcEܵnr_Bߴ�/_j&`��>��M{���'�y��-H��>��"+o�>�,�T@�OؕP�� �Ư�Z�O���'�lr+�A�n6K�Z
q��Z����Y2�w���tv��k��h��⁋g�7�5/�y�R4�����CvG���g��q��
��Ss��B��
�QЉ�-3�R}d@��ra�iA��'��uQ �W�`��ğ�����~����Rt�a���Q��f���c�0֭, _�Ɗ@gSg7�r,�~b���p\�}��M~�/�� �ze�0$Q^~Cv�oK�|!A;�{>ի �e�p������}�8�fP�ل��]���7	��.��zMi���!ipש�z�6�yU0�h�����R�*~�l0������3�]�5����]-�ݏ�����}�˴��P�k�ϡ��렩+^oQN ���	+�����~<̦�6���c�Q�n�}�s�S�]+z����~��s[�OG�Y��¢.��iI9s���nA�%Z˵ϱ�ƒ�ln`����*�6��+�N5�̷D��t����X����2;�af����<cKk
����	�jt�}��]S�Hv���t�y�wt=o�x�Yw@=���8�瓂��/���
���5ޕ�y(}�HĊ����l�^���5ȅ�߫��\�گ{���(;9���SN�i�;#��¤��S#J��Lf�\o:%���J}���8��ri���";�X2g��l:��u��܉�9�2�6����1��憺/����i&w�ZiS�k�֔/�My'�=���av��'�B��h>��"��--���K���;(w�w7�r�����u}��K��/���pW�b��X#1�F&l�_���*B�,���Rm.����,!��G<�F���A���O��{Y������ZE~od�XC!��ŧ-����r�?k�_���	V�I7��� ����6�]�AN�)�r9O��%�&t� x{թ='�/W��h���L,�}��X��B�#f���i%�Z�ޝ.�w]Cq�p&MϧKm����u.�rZ�^:7�����)�G�Kt	�C'�MW��ʉ[���Iv�k�����tA�:E]���ې@�N@'W�����ܸ��z/u̡ν��qQ7��s���.l�	f(�����t�+nW�2�]���C���|�_d�|�O޽�G��#�O�Tz6(R��RjI���!�D�z&,�,xtw!�|���9�,�ȏ��.nk{$���L�Đ�D{���z��k@L����f���wݖ���,�q֏?��s�am�.6D��ݜ���c��r4ծÐ܌�-�d��7r��a���.m��W�_��b��QhN�7dMqe��F�vE.��8�~Ww��O�ӻzp���ZP�i�.�������.��h7��/�;.�fn����A��T;d�|�ݳ��)wP3ܰV��)��]��a���{�!���h��Rռ8<(p�|��܁}	��Kd@t��� ���%��!���o[�inv4 z��u��rO|�$����f�.�"]:�6�|�Ϟ�&�J�`���T�C�CTq ��2��>� �~���`T��4)��DNZ�9�O�}�LZ��)�O����`�{[�ri3�Y�M>^^��L}����j�Z}�dg�Q�+�4�=�5[��(do"���^�R5yV��QJ�d�)�����u&*������dϝTزg�2K��-g�Qnw
@�����ύ��Wr9����C�񕓃5�}����Rv��\�t�i���@�-=�J�l�I�CA�*��߭WaG�u�p�Z#3D��R7¨o�I�q����4. g��+WwT=L���$��t��z��{���\�� >� a���r����b�7jp�hw^XK�����9@+unj��c�U\� ��-��q�'aB�^>��v] [�5��5΅ש�[����g9����2�;�y���8][g(�"^0��3."�:��k�m3����������!�(aS8��SZP�g���+��JD���'>Q|-�,������ `b@ת��#n ;*��2y��x
o�^�QP�!Ť�f�n<sG�_͆���13�@C4�K��8�KaV0�Ώ��ə��TG�94`�bN�E��>!�MlF��j{lD�7�xOn���!I�rw-/����er���x�IWxX[\0|�#���u1n5b�{�@&��O+�t��y�c/ �6X��c�����)!d�+�8ϓVOۑM��<��Q7�h��B]�'v�e��������Zl�f��������K����9Weq�A�@ă3�����Ԓ������q��)���Xe*��jN玷�����ntء8>-w�[d·�5������?���� l���!$`F9W�ˠ��zRA�������2�gC�yhW^Ip�	�B+�����$��%����$g^0B˨�S�nM�!x��p�`�Er�4�1�>�����^`�npq�i��c�H�� ��.e�6���
��Z� Ӣ��x�	$ |2F�1�O7�]�ܖ���˝җY.p<.�_��������Ng�z�	t��jӗ&&�ixzf��� #��+	T�-U����hs�2e�'g/x��c�9s��^�U՗a��X4q���h��Qh�i�Z'����0[������C{[�(�1cG_z��u�/`��R^��i\�wP�'a6˶7x�S.Y������~��5Է4ʔq��Ov01�Q�3���g5a{ﺣc�4�k:��*���m1�3�aӌ�܂q\��H-A~��i4ݺZ�z�q8b�p&�	���K4���FH� ��k�V�?$Q�|^��,흚���F��I�b��'h�2��'������fĩ.i_G�!��<{�Z4��c��ͅg�#�Z�H���Cb?w�.��흏���s��fE��a*�kf%���C��mɸ8]	g�;���]h�%i���1��H�T���1a��� �d�Y�cJן����v�G�-;��v׽����?p�,;�u�"'�7�!�<���g�D�ƺ6��g;M�VM�3�䅚R�������}`��%%�pY(���q�@0�{@�
$�D�x75*�N7Σ!��s���N���,6ր���rb�=�"�Z���˼8�������K�<l�2&|�.g6|��-�ǳ@��8y,�7��H^W�H|t��!����6��q�z�ō15��:�ݾ���T���A?g%EK��.��ٺ�z"��Cq��7ܞ�+�2��(��^JXsh��7F X��� ]XoʊOފ��Wd4h��0M��`#o_V���l�����⩐8���0K��a�B�wVϧ���m ���g^���[*����ub�H~E�%�`�.�-ߝ#ie�1���>����A�#(��h���0F:����]V{Z�5�f��u��3���rjA�!��Fp��n���!�i�B��y�b)�6-����(�:t�_�Z��zu��%��X��Ĭ�B�U���d��<[:�nz��&E�����aD���L�>a��۔R-��qPa���5[f���I�
5�xA����P��Dާ�0*ɤ\��o�f�X����	}ͳ��齝a�XZ�v����v�^�y�*Дʹ�����/�H
Q������5�I0(f_��N��0��dG�ҒR�c�}Z��b��䀟�t�W6d&���7$9e%��s��{��8>K�j�:�l��K�["�Q��f��⚂|�<��W'���H7�޴�l#'D&O��\��_M����El���y��L��TB�"��dHwxlj�7�i�����ќ#�!�����hb�8���[w����dp��ʃ��so��,ߛ����Nf��O�S�d�Z��s�^�����QGG���O�I���I����%Oe���z�k�0�z<\X ��6UK,KLh��(&Eyy�ִ��>2���^�2v�L+�V��a��jv����M�k�>����y�Jt֢ֆ�l��41�Z?��.��ٱ��;�!��&+�����ʪw�;V`�D�@����#q��zU���t�c��ܲ�D�F��9af%��M�R��k�9������?dh;�ï�h�(*$kP���W�o�T �>]d�P̏�e*ز-�9�e5�7����ջ����_��5�q7;��Tw����4�*3Њ��A��Vi�Y�{��Uv	�G�:`�3�.Lk�W%R�]xn�];V�ZE����k��ƧN�r]�:�Ah>�����)	�vj�`ݙ�"�a�5P�t��C�;,�z��t��J�f�k��-q�T��*ـb�Z�s��7�w�{K|F|bѼ�~�ڳKY?́ںdd�\�f@u�بj��R���N(��u