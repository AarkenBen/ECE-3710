XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���EH�$03n�K�9�� ����N�W�k�FwO3*t5�3���K�K�kA�N'�'E���U�r��\���
}�� 8�����Ot:�-���<��P ���O�oQ,D�..��0�(�@��֥ ��uƘ�xq*���h��0�;��}����r܌�����a!�	��y��)�@ҽ�����$�UV�t��+�-
����m_w�4���� ܙh�"Rzc�/�҈�zE�Wp�����~i���W9�|>�Ah�諪M��j.�}�9�3�t�`$�x�q�֙���)����t�5aA���(��͛
� ]�]f	~�T��{2���,J3��_��i	�~,r�V�M6�H?�t+b���S���Ms�T���_�G�A>+� ̕�4�T.68[���yr>&i�.zz��#d#6�Yŭ8��i�����/2�#��x�����£N� �v8��*'����� ��z4�a!��RX�sͮd��'����)���S@"!f
5^D��U��e�݆6�2α_�k�O�.L����iO��ꥮ���'��*�)PW(��s:$6o��8��R
�Y�c��^��[�Z_os9M@A����J���;�p�{���K��Hh����V�fÖl���-t��@S<-��a~Z2HP�5C;�9ق%�ǘ>!f�%� ��x�[�����^@2Qeŷ�&��ixqHx~�	�Z��AX(@�\B�*�[�T���?"�	�� �m��
XlxVHYEB    b8a6    1ac0j����P��DB��pl ���B}Ǥ�0��s�a(���)��,U���*ߧ�Rr�<X��-17�˻����gA����J�n�ĝ����ˊ�^��tA5nn�8�w�� �5���Dq��pЄ���>�i��7CY�C�?(��U�Hr�=��h���:^�d��J`۵� ���-�Dc��
�:Nk2��*�tȝ$�]�e���o5�c/Z� ��A��)�3�XwP���͝��b�}���;x=O '�儂�Mo%�h��ԩ�a8c���A��Ϝ�4�Q! ���0���������Um"ɧ�Q9u�x߻X	������-�d�}3Mm��y3*�x�Q�F���u�K�1
���G��zi��f�50���m)�O�����<�CI�nffi��d���^a�r�v��˼�.C�������C�Pv��ᏆFaWH��5͌\NZ��BF�� Dp� ������U��4u^��R"��AY�i�����nb�'߳V~(*6X�)����������;��m�%Gr����ܩ�:�0*>H����a�{ǯ��A�_�����o�_}�L �3gI��kEI��938 u(�^�fu�8�8����y�u���[��R����A�'V�����j���Sҕ):���'C��W`�ab��ڝ���n@�ru�`��!B;v�^���S�jΐCJ ������@����܄@\/�;VO�h�"Ui�r�3�艖zi�)������ےO
)���S�9�n9�N�';�Rm�8�=S�X3u�7$���r�xN8�c�b���)�8Uғ�G�w�c��>|��)�O�,}_���6Z5��('��D��a�܊$�{��!5[�vO�{ʌ:�����B~?��p�Q&�Y��d뒫b3���D4&�Բ�{7e	� �Df�_�����oJ�~���x�!9e�)�{&4�\�@X����aƐ%��C�s9-φ���E��w�KV�\B�n�Y�ix^�����q~1?�j�����.Ǵ�O�f'�z����p�_%l��k^=9�]{9�pm�	&��ٗ�w��^��y��R�E9�P}��[�!I*a��)�Ƨ�NGys��T�X���I��5i$�9��hqdgB�u����M|�S�ga��љ#"g����і~���3}횒p���,yb�"�ʷnK���oL���K��f+I�r��������'E�9�2m�-�ó,XC�B��b�#*�#\⨮�䕾����<>dH���o�A�j���=#�>�uuyĊV�����U[�'�*w� ���?>`[i:�e����T"ᜪ|o���쑆F��nR�;��3m穝$� q�l���C�{� ��h�r'�p�]w
l����B���6�f�j$9�n����l�T����K��z�*ZN~d�k;g-j��C($L��gl4Q�V�c�sP��Y�Y�?��W�D���@)u��X����B���+�)}赪�Y�Βr��)���ݛ�w%PM���*�84Y�$���g!e��g���F#�)����ٹ�)�fDٷ�_��Q�$�U�M3���Z*�ֹ�{RQ�kR��vX���s�tE�<td͚�ixh���C�/�J�B��?�l�&�w�Rʉ�
N��.�l��t�|����p<s�5�ARR�h��9W�<C�jr'����W[�o:5�����MH5�Ց0�/��g8WI��xّ��CF�B���\ή/��������ۭ1(`LJ���?����Yb~��|�]�����X�{�����!M������'R��PJ������� ,?դf���*��Z_�6e܋��s���
���Fm1ה~�K�h��Т�?aD�o?� �
�-;ؾ�B����΃�GtSI�Ir� �	 �j�]u�P�1���p$~��S�<Bq[$O��#�[�`�?=����J�.�;��P��U~�����͸1���95�,�J��}�$ʣ�.Ƿ�8��0�-l��3����!J[t�4S7$y�'���`UH2�i���	�\��Lv*����KΚ.�)7R��>�RS5(�ɬ˳��F���[��n&���Uq  F�<�|��#�T�����0�f����Gj��p��WԿA���G`�%��s#��2V#�����B9>n�leٳ�$�5q�w;��>� ��+^H���z�.�_�<:)�}o�y�Gnoݭ1ĲΘlOxf�����[Y<�0BM��aYHή�A��D����&�u2�����u�.�R�r�_%�zJ�n��7�F�cEp�h��12�a6�t��~�����,��=	y�U�����؁����P��s�e�bR.��w��Ċ�#Zs|��=���rҒ�NlvL 50�_ `&��_[���*�E,Q��R�.bT����O��90���ȧ���5x�H�h�xG���x�(8�<�m!*��#�aʠ��C(I�m��Ag�b8�w� A�꾧�i��ej�J�$�\�ivs5�w��<�����T��V!�Z�I,��i@��&鶿M��V���*���c�TDJ�֏�>M��Qn�������
�(y��x�"н�����ك��Ŕ���M�}��/Y�+�E�zE���w�y��_�sF�ٝ>�wh�Zi��q��<N<��ԁt}#r�pSm�$O�/oWED(j�T�M8�饽M�K[��o��~N$T�Fcl�&.&3�!�>��t7��;��cC��a�%}��
����|�k۪�8ȽuU�םzئ��0vJ���,^01_L����n��(�*9kc������]������-$unn?1A�p���	���≀���X�����T�@��(_,�H{Gx�SP�H{y��W��;�jN���W:@~�,Z����9���q�
�[!+eb��*���ݒ&�e���h��ܦ{^���uNS��K�EM����{s���q�7A	�h48�����r��"��7+ ��F����:� ��(�4�&w߼�|V_	>�1�̙S�[X>R��b��	$9n�C*��qGJ���)������<�(�iZQHQ�B�
���c���j�S�&CǢ=�?��ަ�Kn�:ql ���s˩�ʰM���0�M���{o]7bS��7�1�g��F��1�;�6v`;g�}U{:��"?��|/�`i؏��D� �D4�P~ʗ�z|��(�ۑ���Cd�XmT��%pgf�nǀ�0�=xSԶP쩸���C1����i 0�j���i��B�`�LFM����x)x�lW��O���g&��0���Z��:C�=���z`�;^�ki5'���	��U# ��T�nmb��gG����{��<PI����M�(?<t��<�(��Pk«e���ի�5h,�I��5<N���d�����xV]"�W���7�z50�F\�1�
`�i� �-[��As��8 K���.U|ac�Pڻ�9w'?q�F�xX�n����b��N�� Q����cEZ,�yx�cּK���u�g�s��Ez����Ս�^�bE\o����S�?u�����S�?��A�]MJ�X���x<��������{ ������<g��*}�K�d#�
���Z���Ͽco9�� �;�H֢����E����n(�Hۛ<f��r��DLgƉ&Z��gM���m��<-�;r:�����qA|mܼ�L}હ8�_���K�j0rG��5�Kc
f�`8��&k*��.��K�R�'֖:��w���q��b��*b��SҮ]Q�H����$s����w��P���Đ�Q�ާW������Z��>[+�N�:���Z,��������(�����h;M��\�ؘ��F��\��^�;Eg�y��6}/nY r�p�|����������#��Z~iw|�E��\�5�}����p}�u����MBaڭ��(��|j�Ր��~^����fF𶳚��%�-�9o~kN�~p���8�!�*���͒b����?�R>���;^�5F6��� �l�XZ��GBȀ���t��Ww.-��*��¼\���k�IA�l3ReN�s��0��`��>��sUg_�2z��4�e�va��Ep�F�P��.����<���)r^���#��6���$���	�&���"�:b������`M�FU��v�FM/����<�h��(���ȟ{�������h���O�:�nx>�ZMk���ח�[#	�\�!$:o��*�����:�{��h>:�=z�GW�{`zIΕ����e��X� J��O¯�ؔ����xҗ��9���7u,_���i��9S��^���5U�#Z�hKX����L���y�Ex��u��>�����[���.9��eĕeNES��CA�w6n ���	������}���O����G4�sN�RH�Y�u��:��q޳^O�]P�n����;8�~{M���\_m�B>uJWO�	:�K�p����� /�vz��2����Rx��� F��N��VTۤm���>����J^�=�}����3����ڃCXa���T��>����j|o�g!H`�b�S(������*�+.�$g� �E���ڮ�c�J�������v���4�QFth����n���9d��~ٛ�.���q^G�X�=G[���C�\tJaK�����JUV�C�{!�-2]��N�@bꉳ��\�4h��z�/�R}!�B��,�����<c���;�(�P�І������
�D�_�';YUb5pG�I�H!&�5˾W���s�]fP��׹�?��}���2��@�JTW��f�u�g�������Y3 bj����l�2c*6G=av~h�1���h��2,�ew���(������5S\��3�'�Q��6JA���	D���G�� ����hyں �b�`h�t�b��en��I����l�"�r/R�AMm�΄d|(#ly7����b��8��"���E�ޅq>^�c��|�V�H�%�(��
-��v�1қa�*�Տ���4����a0=h��Ṏ�D�|mƾ5뉭`'�%�A2����R�X�I�]w*��h�e{Ầao|�	#�5*{�1� ���t�i]����Ŕ�/	�龬A[-6��I�S�h�)�c�����G�갛B�1Y�j�~�%�5�bj1�����'6�WDM9�c�>�y�F�M���|�������ʋ����¡���m�"J��� \c|)ˤZ)D5w��t�C	���d���	��)��L�G����ߓ�� ��+9j܌�ty�ɫɝA���+HwUN��kxg�(�#fdrS�c��sB��6�+�0=��A������p�u*+�>��`��J��ߞ�A���`��G�ʿA �C���\�!'��/�̺~ּ2����.����2�f<�9���4؟�p�P�����@a*�n��l����Z^{V������a¥ۘ��s��#�+%�*��o�gd���2~����$ݭ�g/q[�<��k�ؤ��Q���N�,������~��_�#5�hvY,R����CY9����@/�v��6��ʵ��>r�X�I�~��q�.`Q�O�Àz��g�Q�p ؜��[hƻ����y��3�Er	�v??x���r 2�c�A��[�k�W�����4^�T�ۏ�qE����iD��kK��-��],���Z��Pm���4���[�ߔ�K*
����tV�_���|�G&��찹�0-�K��SE��PV��[*��	ܨȜg��#��L�<a��h�W�J���ʮc�	�0^;��{�w ���2_���)��~��/�^�w�����r��}I�
.4\��Zi$K�����m!�"�5VEk��}�b��A�
���9q��Vٕmw����Yi[�"
x�ƽ�Q�v鍠"�����l6<�W�z5G�I�? ��O����U�@�� t����sJ��`�~�>�(I�tj�n���մ���~����6�|j3n�]*�2!��j���7rUj��48�Q���TM�~��_�SkW�z��)}8v�FG�/~!	h�{��b�S�	�M�Z/T���-��.0�s�f�|���NV���۟�OK弬�JL��vi�/]{�z�;3P,�Qک�'�:�>]Sd���P�A�'&���S/�$K!6,+�'��82��4��%]��A�_�����"e"L�<=m�ru�:�M�4�'] �`5u����,���=˅v��	`䇱_�����$��"繩���7z�p�;ҩxyNY"��y��"~��*���V�=	����	Rv3����}��[�~}�޵R?�u��b�a���_�F.ҰӼ9ҧ����b\��/��l��ͫ�L���7A���;�tk鐨�o6��VG���������E�4�W^������i ����k�0(7ױߞ���b}U�+(_�*����zP|5�l.�;�_�ڟs�e��r_Y9*��K��q5����u�n"�&��9��l}��lw�i���FN�	^�;��x��4Ka�(�_���PE���]��˪ݚ���G��{/���]v�9P�Ko�������`Tï��BOO��6��!`��Q�W]`ȣB���v@�8�O�:�]���g��b?��?Fz���z�]|��6T���)1|����m�x�+�rP"f����� �d��ǓU�7E�^ҏn]�/(�3�z���B&��.�4�Z? �s�����R&