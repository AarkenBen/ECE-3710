XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C\2���WtO�����-u�:@&h�L������`OA���g��񭗂M�N�U$\2����p%�D[���}�x?x/�8A/]r�*��].�c�w ��͡0�����Ğ��ia�
���Vyu2! ��B@ ��q:��(<[I��@�M�GY�)r1�uA%�yg.]���!;:2���h�?�j����S�|^��ld���&��82g���b�I\y�ڀe8�@��#Ƚ�˙(zU�����[y��@���L��G��$UGo��FA�&{���6����)ɭ�p�)r��j���[�pat
W�a5i9?U�_��4#؀By�@�9�;��B0��gU�&[˃м%F��G�Ϻ�X��7Pŗ��	f��D1�;�G��@y}rr�I�	�Wݡ6˜�0�y�y��@R����b�<���|�����{6�������`�ce�G3@ω`_c���j;o���*�u&t�*�P+�,L�O��TJ4��B幕��J�ol3���2���[���b� x7�z���g�Q�@�+j�P齮�\陌� ��ظ���]\.�ꤚ����}��a�~7���q����9a�c`�Ԇ��݃�q��nf0١I 2����2�$ ��7�����=����X�K�Hg��C�����s({��q^�P���]�j
.�]Z��]��)��Hܕ���v�֋�Azi%V�C��a��
F&�!v��=��g�uY�����OߣD����XlxVHYEB    2e55     b00@�5��C##���E��雀X:�����2Q����\Y���bh����v�������?򅠽��̯Cs�%C
���8�8�j!)�����#A�Y<�ל��G�Q����J)I�oy�J>�T@au�(�C���6��������{�c͞� �%�z�(zV�|l9���IS�5HϤ��~Ha�W:���uB�J����/�cFU�	��=���"#�!�@�T��PΩKQ���jt�O[%!8�W��Y��ƽ�78v�����6�h�%[?na��0��0GM����#f���`��&Y�8\ԋ[�rs�/�>�߿�'Q!�(�C{�B|������3���ӱ}J���cM�Č��� ca*�m��hKbq����e�е���H��]l�XJ���D��[��J՝}�o���u�����C�fGĎ~,�� &9�X������e�)�H�)n�& ���[Kا\�`�"q�L�|S&ZyJ�w��Y)�UÒu}���o�t�I]�A���-|N����\r�k��{��t�����ݿ_�g�u���pJ��ohX/ikw�y�AS�~36w��� �XW��EvS�������Y�ι�I�x���n�h�v�7��S��F"܃(�K%�)�r�P%��a�܍�K�Q!����hTI,�L�S�HR}�:��o!eL�ѹ_@�0À`���իk^G튮^1�%"�{�Y�A���G�T�@�t�:bj/�
Dn�����7]Y8)ߔ=:�;���b����%�z8���}�)/�ot�b���7Ĵ����]�JF4�Nf�ZGy����6��3���ޔs�[��f$n�U2�����4�H�#fg#��p������>����o��)�n��D�^�A��q�{}�[QL�A���C���![iѾ������ݣ�|�^s0��J�&pĈg��Xp�"0��U&�^���x1�U@��hd��[zr�$He�UA�R+U����gށ�Q��M�4�6F���8���C<�r��1T�	�vf��\
���3�"�E�I��f�WOH�Y|�ܵ~j�����6P+Vi�����[l�.�S���V��E(DB|������|>��9���~H�F�j�l��,��9/ǂu_�>_O�S�jc��'�~;�24� ���Y�th�x�����<O7��({mS�[QV^/d?��i�N�h�����|�i$@N�P�ᮗC���'o�����!ۍۻs?H�-�9̦�� 2I$�9��b�Wc�q�S����1)/�����3DSb�����V�����*0�%�G\�3�쾒���𐣬XXz�Ž�<�����`HN�i��|�_av4��w�% ���L3X$̥�m��W��K�۰Y�)��'B4�@�;�}�31��2/�'vb#M���������6�����|A���i4��D9,��X�A�c΄
C���G��d�V�'��~�[���6G��G�#}bl�<
^t��-���dF9�FR�G�J�����J3N#�Z�aqߦ| 1C��GǍg!�\q��g�����k]j��4�{f�_�M��4iN%^W�B���{9���>�P+�k����S؏դ6���I�\I��[4e
��H���o���t�H���\
Y�TH �X�����<�v�"��a�FB�!'5*�Bm@I��]�T<S{a�_��ɾ���4��k*���=���\ꕬ�+-�럱��bY�Zsҩޥ�"�jT�?���1�(_Y���9f�Ac^s�a8��o��7(�tפ�^1䈏Y�n�%3��j$�Sv|l������]yR�o��s}�_'D
��D���6�pxY/��y������urB�m�����D\z�{[�N����t�vͯ 	�-���x�tCZ���&xb�XAm�*�h��û}(0���i4V/� ���}���:� �n��0�.} �I�H�Ҍ�lrӰ�u<�ћ�$[ �*��M}��c�(�j1ΩB�گ\����ē�3o��
���"�����c^��y���W80�E�ٌ �-$�|�����������Q���Y]��������d��,��æo��m��O/�ǎHomx?��l"����O��r$��Ą��&U���ui���A��P�l����{��[�s��1��0D��6#��S/�BT���-�v��
 �w�+/w؉���t;m`�s����y�3bI��j�p��8hh�44(@�	�g?�&^xB
��6�[�����F|Ԯ�QH}��΋��\"���`۠?���9AU��:xR*z���3��A�|~��AHc�7=*}{�ڒ!@����hG�#nv?j�K���S�Q* #�^�퓅�ff�
��f�KeTҪ!��U�L#tc2�考��4)uL3x��[��y�v�hIҾ3���L������!w�b��A�D���E	����{�a�46�?������"k��m��D�gR�{�������3��u�]�ط�f��˩�K��.��><��h�U�F�aIve'�a��/�QpÄF�:)A�3�T;.P�Z���P	:�*r��i�D�����畝�y�[Xk�'��jG�F�Մ�r��x�QY��pXLU�j{��w�
�O3�����Ǧz)�w=���n��W+Q��3��4>��z�H��F�a��}ޢ.�7�~Y����6̪~�3�@��a�m��5_bd�c�$�R|�m2��'%O6�ޛ�c��+�'����q��ǉ�4���=w�I�=��_�