XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ޡޮ��rv�}d�{��VO3yD�S!	�d��:Hv�5Ɣ+����6��b��v5�+��C����H�_s���Ӷ�����h�%]��H ޕ�!��b�g�?H�x(2�i>������хs�ӻ(=��5Dr0�uL�5L�
��l�=�v�bo"I�m+�|az�,
�J�ξ����������g��嵪�s*LjZ�vT�cL��	�Z�Q9Y"�2H>�� ��o]ے� �ಛE8��"������Jx�1&�Tە�@:�����hE���As�u�q��4<�c���g�U����F��:pl��ឰ��/f%�KU��X6�:�1��:��$���g�%��L ���kU��7�X�(�MCV�.�b�m�x'g�l$@����= ��vĜmu�~�\����Si����Hd�ľ��r�!�<��N���*��(�zm�*��`�&�os#`R�0ĔP�7���E��TK��e�<� ���둣F@��yaGܬ�EJn:�QW�Eα�,�9�D	�~�]}p�	,K��?'혨���]��I���5�-�_�	����ж��o8A����"���`�~�c��ˌ��Zxut����0���Ly��0�U�Ȱ������#|��k�V��v��-dJ���Z��!����lv�e�PJF$�u����ʐ��x4,�-�4�ڇ��!�;y>"A=����W�^�rpţ�5ء:�
�� hb�iҌfV0YORYew��n 1rw>مj���gk1�?{�CcKa�.@x�F{��XlxVHYEB    b8a6    1ac0��	�3����jnvj~$9\� ci�IG �ccoqnm
;{�����!?݃&-h�],�� �F���6x���*�c���Ae���?6f<BU��m���N�kҍ��S� �rߋ�6�:���\]$*�?�
�Ϣ!�"EJ$��Ȯ��̧E���Df�?��Q�RL��N��e�U���#��l�����ՓuG4sr[Z���ipnn������|��hRx�Fr=� ������@�K��m�֙�b�#~�����DD��R�u�A_�͑.���͞;��㝮��M��Dmd�Z�qK�ㄍt��и/p_W��羒�'{Q�(�p/J�v+K����$�t��tg���-I�D8��j% |�$�m9.��}no�=�k7��r���gw��wz�F쎑��寒+\����r�pʢF��:,J���;�SFHa-���B�5�G��;�!T��Pk@�gH�����]�R_�J�x�y2�n@�ڨ)��Wk`@��,��������"�ۋ�Z�{�s���.������T9파��gSM�Z(�݇�272��-h!��um��~�3���R=�3-��>���Z����>��H���B��F���;��8���Q��&�3/soT�(0	8(��鶱'�&m�}(d
��_�Y�����Tb�6�l�)��I�����4I��m�qDQ�̭�����
�jf-�J!�� ��<P�W��]X���hj�|�C��]����-~Z���t&ȑmt�mZ� ��p�� �ܵc�`Y;WA*!Q��K���*^&�7��5�;3��Wޞ�_~APX�%������Y���RB4ae��	�c�w-!��א��t�1����ofĐ�A�
 �wۼ�2VS�=�����R����;|�m8O������~Q �C�@�_�vI5��ڳ$�aړ�Cs�B�dQ��7�Z��)��'���"m׉�9& �  �N�4>�N-�+`���f���@�0��N��7���s  ҒJ�h�z1�*�a�RL
���F�yN� �/����YVi�T�N{^��'�J�vb�ۿtJ�^�u�{��Ǆ���7����[�m�LY�JjK��ʊ���f�/��w��Hc�����9P'U�{�Oepd���|p���j���-ߡ�w���V)$&�]�ݍ��Om��Ѣ��FT�{C�v��a8�؄�>�U�xm㼦a�lw����EN���k1��SH�q,�O�\�Yu�TBR5��z��ʍiϗ�������d~aU8��l4��f�$�E�"��V�n,��.�~wB�r� {�T���:�����x�[U����u.����� �e� ��sC�N��:#��\=�'��(�����!R�J*SQ�RvE+�3�5ڈ��8X��x�c�o�
Q��A��Ї����[����w�˸YH�l�O)�Oi�?b�?��L��|nY�'�MʱYz~	��`䵾��a;!e�ʞ�����[|� V2W�Q�Bhz��~6k�E����l
L�]�ӢF�;���ۮP�7!����[#$�UH�4��!ڜ�[��|T��*j}T��V#���s8$*����*�����m�������a4x$Y2m~a���\7p]4̒���R�'��o���}8�7�����>�b��h�Y�9��5��K{#ވ��҂��!�c�u���3;Q�c�i�FW����QT�4�^'�%?ٵ�Z܊�HQF�Nm��([⾧������		�k�������ω TFY]�J��r��e A�m4��21�k0{X�M�����钘�?�H�h�^F$��g��؅�~��..�,�9��XMltCQ�ʨ2���)��Gcғ7���Jb��$�k3��3S�qG��8��_GFQ�ۈ-����y��w5)�J%��H�I�y|�N���� ��o�K��"��7��+�x�PA�; M��Nn�I�)Y�y�i�Q��y��ta{y��/��,z8�-4�{įRZ�	��VN�8a3y|�a��Қ#���V���5���C��S�FPt���Ƚ�}zMz�k���]��|��:�?��]�ʤj_,d��f��ۉة�A`6���wG�:8��
"g&m��5,�ˠ�EMp�z�N�w~]��BU�b��wCVh
�&�	i��VJ��7p�IU7���A�����ݾ��D~n���-M[X%I��-�[�����(�V�Ka��Z��5��Q��)�T[�O�i�q���O�7��1Ƒm��Y�g��Tً����z�<�n6��3F
��!oZ�bz�o��ߠ�Y`"���çiJy+������	��L�j�7�V�@f�Q!��ܮ��v���#�ߙ�1��Q�E�@{�^u��O����>�x����'�HV��s�`�l���:$]G�(ynm���6 �"&�Mh��Q��CX��O�S���-ɂ<D���k^��Ṗ��	H�1.���@�#��u.����W�!�o�r� ; r�%�1+x�We���f�[\k��R��7�	>k�/'�����۞w���/D]"c�Y��c, �WuԿg2!_�K��9x�U	���fuŪ�g�T��{xr]P��?�e�R��tZ���L?|�06?P՞C)~3������g֘J���EH��ѱ7��a=͇�;�����;�#���c3'���=z��{��P���N ��j
��i���o��Kڙ%��:�������%/�|�	[�^���9��@t�2}�'�!��ߛ������2_G>f=:��Ȥ�w�<��m<F�߰1��ۑ�p��J&X7�l�����(e���o���S������{�g<�Exh���W%���9��EyӋSB�>')L��m��Lt���l����^H���I�r��Ђ��!?�|Ƃ�2�/M��,QaQ!e|�-��s��~���˒���;�����@�:_�C����Ks�u��h��I�[��u����}Z�P����[�3!p�H�S9�7�|���]�5�����]>�P.o1��Jc�Q�����c�)X|�]�[�F�/$�(]�QO4���旒O?�Ct���N\�;Ys�:���s�����? 2-�*b�6��P�n�V��Q��`�V�*U��������m�xj��t�� �>��8�	�� ����1t�Ń�Li�wr�;��,ƁMiGv���S~�CbKZ0�k�\�������z��jz㊐�X�Pp�`��?Ea҇�^5����9౞�g��L�K�`I�����<`B6�(9��7��2k�H��R�RH��:	�Ԭ�*�[*Ƌ�W���2�gz0�*�❺"���E� � `RVX��I"p��= ���B<���'�r��;Ys'��H��R����0��2Ǩ魄�/^p������U��?G�	L�;yxᪧ/��_�IM�lsn/�JF�j����q���B��랐pTS�cׇ�1���gq��p�;v���C��\M4⇹�7�6~�|@0Y�^�&��h~����j���5��T��-��۪a�R,�X����`ol_dMc>�N&w,�j��,�|�y����@������*�!�(աn�+�C;`����M�� Y���oT�S*By��g�ܞ"��S����3�޴�G3�^M.��K��4t�+0����ᝋ�hj̼���Ļ��6_��H���-�0
�2?C��|S���%,t�@L��N�K�l�8�W��B6���X��Ζ�5�`�K�{X+�e_n�����p��ث$U�{��qQ��=�	Q"�W`_>�*
��E9�!�y�H���u5<�(?��ėZ&���[9�ă!zw�kg�0�����`!���nn$�X啄�{k{�3��%�٧y�l#���#	%K� ӱ+��鶸�w�x+��W��Ac_�#�5Z�!ѕǡRAG�tK}���=)6�Wb�&a�v�FkA8���n�<]� x��-��"z98�B����j���8ڛ�4� �0��v�
�%u��$�3��UGe��З'M8{��g�
vu��s%�+��vk���!���k<`�3��Q���,0I��5��;ly��*��jX@)a�sՀ ��O�xa�ytYg������.v%�RT����x�}���$�baE���%�dj!0�uW\ĢI�+��/�X/1éP.�_|N4�}+����_��n�z��b�P�&�u{���rx��<���$d���� 6c&��̽Cf��S_�0�FL�h�ȲsE�bY�d�^�^Z���޲�*_.*7j�c���G�H��ܹ����a�^vP���w!�8���/��G� ��cە�֛��m˕�eAb�Vh��En�ї�_ɱ����NdH᤽�@U���Y㽨�0���)�����t���f1��"W�u]����kM�Ʊ~R��,���z�l�Ec�\��ʱZexN�J;'��Ƽҫ���+�
N�u%�8ѧ��a�f�R
���"�Ǎ�,-���5OS�d/ �i��8O_���O�T�=q)>�)Æ�^�����A_���@��5�g瓺�6`����q6r��-s��Q��em��8��w|M7j'33n�.�������O���A���Kb1	˜BՎ�Ŵ���9�a�q���a�7r��Po�!�\�[i.di1;��{������A9Y�p�i���%���@�|��ݕz�s��ݤ߇=��lBy�ے˥�	�=�n���L�B9G5Y��f�/�����f�7N�����C�L\��p(��u�߳��z�%Vz�;`��c$�S�Z\��ȕ�zo�q��0༐4fB���9H�N���_����5S���8ￗ���i��i�����S�
�����w���Zm�̆�.-��i ÷:+�bk�����{���G��zcS�?���1�*sh�ᐜ�����\��Y�����t�gG@erI;�������^FԘG?L�5=h|��@��(�Ƶ�+�*2�qM��H�+qk$��3eH�-tk4q�4Y���]����L�ZS�Q%�H�z�bї���*r\��͸8j��PuC����z���z�ָ��Ƴ.P�5�^	i��vuL��ۇS���Ý�E^�wa�˾<�Zϗ��F�כ�b���H���v>����nNګ�(�9�䄝o4��7ty3�������=_H����ϙ�o�yqL���oV{�-������q)^���'Ԡnbj�	�m��1�׉U��X�	@!w��Q���O6q�7�w���M'��6��	���
������,6�|��h�q�C�M�䝠&~ґ�� A�I�L@����-m@!���­���\:{�gߺX�&�l�v�eo���M#��u�ý0���jl�s�s�f����T�cJ���4(xU�| ^f����J*)%;�,�i�&��wt���!�;�&�ʛ�UE5(
���5�w3�ם��?�V��t�r#��Q�V�o|�)cX�$7{��Sѫv������{�@�F+��U&4MA��k8����1��6d�+��Xd�����O��	�vōϚ6�l+D�v����o�;N/ �%��S�AT�mĞ�����^�9uOơSkqlX��b��+�a�v�P
���~��m����SC�QHL}�`����GH�qT�Ϊ|����I[�����*���U�PB~�@��R�{�$���V����!�l�\�՟�
Z�#�����`�F��h���E�e�;�e�۞�J�	��ժ�Fw��.�JǶn��c�f�R���#r2�a��A������3�yye�U���$K)��E�>�?u]�+g~n
W=�u~(� 6��#�x����6I糁�$s�w�D��܁f��鏃��K�c���b�����L��!)V(,���Y_��C�O�2�9�9�����79h��i�Ck#�4��Hh��N2��1�B�p�R33Y�y�Q�=�N��$lr���=�8���vcá!��GI���CD�~Ɏ���y�G����E���?���%ð{Bg�G┏_�]�ͽ�sA�a,����/�����A*��A�b�^�}m�d��f�r4F6'�I}� �X�C\�v	ӑ.캍�Z��$d�w{��,�Ҙ^�ruއ&�Su�ځ󫚇؄qM]r7NE���� ֫��x�#���&����*������Ȯi�,N�p�N���_�6cˇ�B���(���۰�Aa��K��Q:��D@$��/�~1� ��s�\$^���=�H����Ȏ��,]�g!���e��>��A�a�������k�g�|.��qCא1��v����
8i��4f'��Af�\Bˁʋ�%��3B ҈��F)� h���2j�)A�h �d������y��qj��)�fKeg?L��rY�$�Ih��"p+jE�����:��A��x#~"��0�[J����j6�}��������\�)>`��}9L��q��%Dm!"19b:�����ϵ?�\5��ҏ·+)�OpMXAC�M��t�zr���*\e��O�w ʬ2�Ul���:n��{��o���_��e Gڮ��-�G��¤�q�s<�q����'\+�݅"�{�K�p�f�qJ��H�9�I�e|<puJJ�KM��8D��u���֯*��se�3k�w����L|���
k� ����p���o��.�1t��,�s����6�ؼ㪔�/Hۊ���~���Z?���|W'�