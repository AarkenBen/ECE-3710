XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8nҷEY���S!\��bk/���ye c�3V���'�wj��U�F/���Y�fÃ�ڳ���m�U���:��g��dT�ח�xv`0`O�*������76�B@���?v>�~��
�*���C�W	���1ۑ��Z���n�8��섲����ai�j:vmo�&2&n���O����sܿ]@7OA2��$;�Pu��gM�m=��kH�@����?�g-h�e4 ��v�8�i�bcO�o�b4;�jd~݉�� g�4~� �\�&�Bɏ���9�j�K<��]d��ɉ��?]��N�!����MJ?�I���^�D���49뇩mO�xa�{�p�B�_x3�8UH��$��ǹ��p�l��Ɓd��x
ŧ�/N;5����T� ����Q��O��y�OO��Al�%u�?��}�����W;uG�,�U�4N/p����2(ԙ<��L*�CF�p�7�a�aU�R룰�vh[���&7��Tg��]�@���C̴����~n!z��G��ay����M������O��v����Q�
��߁ǆ쳪������JF�<�A�����q�o�A $�\gh��§�?uZ
�eя�,�D/�}��z�"��z?�Ѫ�G����;b�eZ�[T�o{���l�o�K�z�̴ A&�M^��w{\n�������nBq<���o-���`�el��8Z0B����[��w��W
�u�+�%Rd�0N���5P��ʁ�v1�6ch��{$9�^��bxY�qEр�XlxVHYEB    fa00    2480T�z�Kzq�30OZU���f?�R�5��Z8��ҟ4s֍��Py����^��S<���u�d�v�Ԅ���B�����!���[|0N��
#��T�ԃ��v$GƝ������;q�(��Q}��ϓ�l�W�����e�˭Gy+\��ܬPmd0H>����q�R�7��j�%���������ǒEE���q�_T�/Y8�'�F�:&iVm���qD�L,u_������ً$�eHN��z��+��޷X�u���xm!׳Q��o�Vq�FI�LL4�%uh�8���ZKE�qΏ�Ю(����g�մ|ȗ
mpH�e_��)";�hoG�g�q��U������7����1��<�>��UF/�\ö�(d�&�z���7/b킥�L6��5#�M�f��U�����U�z��_�%���dQi� f�Ĉ�Ѽ	i��H��O2�ӹ��>+v��'
����ض�����ʸcPZ�nx�ԡ'4���� �8Cr�΁|ɜz�g�}�{ш𥘠�4�) y�~�39uw
/7m8�y���x����-���^��d_�w�G|x�� ��(�?K�/�}QZq�u~����h���>�5�N�
��B�=�̜-��u��/� ��������#\(����lId2vj��>v�/To��9��gn�my�h!���A��0ئ�f
�ɑr��v������;6N���M�'�f[����!���Q:�F�}�[[	D� ɨ���n���=�\[4�T��)��'�Px�� ���u}�����-���m���n����` 9�v�\׹>�����Q.<$�O��M��tIu+�"!�m����֐GWV�9�� �9�T������-���?ݱ�z}3���4�!3�W�~��[
���wo;�5ю,�9��XK�����Uڑ�rk�qp*0�*6mh�$\�3%C��?rMEl�tJ��a	=�E��OAy,�w9 	�����:�+_�'J|w����}JD������lA�lm��4��Ş�����$�x������`0���E:u����a0�t�H�t]e�����FغY�J�����Cz`"��t$�?��UR�A'D��![>Q���n\�A�X7�C�jzx}N+݊�b��YP�6�����Ͳ�C��
���۹�%�f3�S�:4/ap��c���:X$�K��=$��-b��� F��ȚJ+��$;-�ts�f����'�21}@jā���F��+S�'˖H:�U�e|�����>LRūi27����|{��K��������AE0��WvK��qT8W�	?t�zM��<�OL�1�6T�����2�����S�](����A�J���z�3:���?�|�cqe�L!��������.x[�V�C,�X_*/ >.l������v���|TR�Wt�r�5�@tL�c^�̢���A����$�K#������b��{q5�Z�`�.!6[���ۊ�����ItD���g$q]F���P�W����.��Rw��v�+]/�c,VI��@1j�=3ITV�T�I�[�nM�w$������1�œ��E�M�56�i5G�;eBpI�����~`Q���t7����Œ|b�1u�����^����C8�-����l4"��)z|p��;�\�"վ?v�!�YH'��S.!q�b����^�%���������>9F������=���"�d���lxt	�`S�xW�3
���w�G
���L���TMf՗�Ѿ��zƻw���֋-ط/�)�����#�5��r>�� Pm�8>6Q�_������p���b<8�L�����uAl��Vq�Q�|Xm�`����G�1�htc��׍���Q�)�c/�f�!6.�T/D��G����a�Q���5���#��b�Na�t>� 9�E
�Zʎ]J��A���׺�औ�;N�)I�d�AV�:���=Z��P�����bfr��W]���Z�2��f�v�r6��D~�ϧ^ʬ!hR��W�0�[F~"(�;d�kM#�DC���rX����#�_0,��!-��؆"A��g�l�c��^�F���4�����$l+0�:s	�[�������T����O��,_�5�M��B$�~IIVE`�2�����;�`t�h��[��N�CcF)�#�s��� �+hd��
d�����;x&hKx��X���#'r0暗���@S��)�͙�G�L�mCC��	��U^�'
�� 0�u�b<h0gD^���'��h�i�������zxm����%�%��U�Ol�e�lv=�+���j+D�[�`S�xs�)E�R�I%+-F�x��!D��^Wlg�gF�I!�0�5�+Tm�S�%�ݳ��`b CMy� �99�*;� �>�nN�]Hд�v\F�\�]e���5H���-7�cO,�����_��<d�x�+��^� ��
2�����G��L����f�q	��-�h���	ڽ�"U`��M�'�M����$]R���"= ��\��]FdU���k����w�˰ 0�m+�%>{A��@��Ɂ��H8��p���X�3�fH�q��A���S j;u�~UY�v&Ԯ�!�x��_@t�`�U��*b�P!�J��*�(���\<o���́#�ǥHH��'��cS�:!�W���r6kfz�b�șu�Y�Qv��O;��j��YG�����Q��ٞc�!"�pW�b�����S�<0�05�zS��+����m�	79�� U8�0D��d+�N���J��
#B�Rb�<)�Kl3n�Q^,ڏY���tsCR �2-��^B)D��vck̿��W\1��Y��5�Y�96V!:���8��~H8�9C��|T0<4�l���.,=2s�$ժ�o��4��=������-��5�"�QYz&eѵT��E�����F��55i��~��J���6�v�T��6�#ȥ7���C�����8����oE��R�M�L��X>hh������}�Xh\���3�e� ��V�0�3��%�u/���cn��}"���$'�w����q�5�P�٪.��$B�-ټ�y��'P��������)��1���1��Q��;�Ú��E0D��v�g��(��HN�2#���cY,�s�3�yxIy�϶U��`��@���I�N����;o���7�I�C��,��nފS�%��N�c�>��L{!=�| >w�:��Yƶk&�e+�/6�lv�P��qG�V &� �>���S=|�?
��k#Z7��~5'"z��]%!�ou�����s���b�5�
Ħ��x��'?pnΌR�޹,˨��]�Lw�P�;>m܋��=�45��]����M����8��,@N-������ЛP�8�##�%[KF?��W2kmz]l>i��/��T�<�-�u�����g)_� ~�D������t2)Q70��f�Q��������\�?�WI,�[����g1�~\|�ܝ�ICb���TQʆ��f�a�2ŝ�����l�+i G�{�
=��_ʙFh�!��9��}*��j�8�c&�$�-���N���r���A�x�^oDu��(d��amX�|�D�h�J���M�%sQ��U���tO�'T�grʜc#�hv�����?K�B�"j�GY�M:qY�Q2GFBw�<����mu�r�ZS8j���{�+ᾙR��O�*?��5x^=S�9�0.�^����{��F��RL5�Yr��O r����~(ʙȨ,ْ6X�wM�B����>����N99��B��`�-(�]9%�&����|Ty�k?����o���ᾰ��$���J�����J�{ӫEHʜ���N���@�J!���(�2���|w�Y�q�nU��G�WT�ڀ���$ʧDk�=z�>�f1�A�o�6����"_j	������Z�C.����]�����&��p��W��~�i{�$$2��#�/ob:\4z�X�$pTa��t$7q���Lt�YKw��vf(�6�C�/��_:�Xa?ϱ��܊ �U�[5<�<tJm�+-}p@w����H�x��fk0�����oIW��t��*����V��Pd�n�C�D�i�櫯��;��0.�Ҳ^��EBk1�x�����*d�ػ���{ r�t�n��x���z�AJ��Eߏ��!�^����\�����F=g��5%r�Fbq��kBv@$�2�I������x��Ӵ뱻=��̈�W�I��5{�e��[�٨������X?���p�.	C���5�.Ewu�ʚL�)O�^�;�{<�;˙\�A�=hw�w�/��S�$�į:��L�L������8v{~!�����yp+&-���У��2�
�|��uY0���|�(���G��܀�sa�0-����N�Dc�/��ҫB��oV����'�x�]�O�o_���qS�;v�#� ��@li"�K�m�C��A�.��(� �rɮ/ �Z�k�R�+W�L�j|^���D����$%�Cqޒǿ�^����#
�3Wߚ d��j�s�7V�u��wG�Ho�놂+7�0�w��H���7���z�Y�9d;H�|w���3P��K���_�5=_�l쪦2:xT��(�sl�Q�93�������
TƿП�y%���wl��Wu�v)��a+U�L^(8$�@�TR͜����8�܎����C�W[��ã���ߒ�YYqB�'���&�?����P���֯�y��{��\���3�*��c�}ׇ9��ywvQR�Vd�����q��6��Y6������}^��2��3 ܧ����SS��ֈ�;t�!����d�V5lг�g�֕R^����o�j7��:eM����<w� "��p�+���ۺ�2�a�����P������*Nl:ٯ� �|F�ۅ3Z}/�I[K�dt�l_�Fy=eaw`����{l��V?�ϕf">�y��G�Oe5��8��1������$Cs���B2a������jOU@	Ic�J��c��?�s>A֚�u��z��/L����c�5Z���c�E�Y�|��)�2����J+��mU�BgK�Q��>8��մ��Xvp|8�D�6~�ީ����9�:s񆚗ˠ>��k_��ۆz�P�lI�k�4�|��-��S�����աz.�r�~P���FT���m�CR����L�)�mH�|���*��t�f��K�l�5�6� sᶾ��.U�v��w�
Ɣ`��u�t��#{���P�8d����-l��#��T�񄶖�����I�N�%�v�N�z�[�*?�ߕd��/��O��Ys�2=;�xl����poYe&l��5 ץ�a�N��n����)4w���#t�1�����b�n}���:f4'1��O�"u(��ns�
�=�lz��yU��E��&L2���2�t�T�M��rE��o�KG7�23�����s�����mj��&���hL��: �1n�3�^!N��K��ݩ!�,Xo/L��k��`��{(�^�v7�SG�X�j1�I�-����:+�]��-0��˽�a>,�j^�h ſ\�6�~.�����s������n�m� ������ޏ\��,�fw���Y_+��L��l��#�.sy�~�:����Jy�t�<k�]�����~a�&�+� �|Y�̋��莲5ՊP�ڐbz�NkѲ7��po��[l����j�Zx;�r&�r�o~L�O��A&�C���f5@Mȥ�*P� 	�5�ҡ����`�#����":���s��
�A|(���a�}�U[.[��[1�f8�3H�����9ZV�*�m�Bǆ�RO��!> ˜(�g������<�u���Q-ȄZ�,�(�j[��w��V�	L
���f��&��Uې����M,��pV&�.	�.=҆<�v�c
Y�gh&��Y"���i@\�Q^������+nY"L�tI�go(tu��7�:���Sq@�`�
�:�����[�1��,14*^?/V�ݩv�ZP��	���0���e�F��u\pEyT�Os�6��O�u;��6hn6�`~p����x�L��
��;p�è[�g�����V�o	ը�w�^ǚb��_�W��H�Ss�����AĆ�2��n�p�L�	Ս�u@^4%]2���J�N�VE��QP����D
��9O���`&B�biN]�Z���;��6M8�:Y%'�y��܇r�{Ԇz��B��{H����F�x^�VCP�"�*źz�j	P%��˞T���6O?"h"[�⳪���B`�%s�Y�!���
�kR�������)���OC�:Ϗz)�eS���'��v�ty�:��(;*�|{�y?��-G�F;M=����h���=�-�M�#���y��_��t+	u/�q��a�W���-& 2�ѓO���O*��$�b���r��R(���1�l��bNK�Ĥ��t�;<�s$X���"*���H�h9�ݧ�01Oy�l����,�����w���0e�o��T�w��3�9|����7&�v8�T偍N���<1��ʎds�����}�5�o5���d5O��en̼�Ճ���R͉�׽~�>��T7��;zv/�Q$�ez���zEB~���%�/h�|�� N�"[s��~Y;������ ��.��V2(���'+e�������ҵ%X`�Y���nU;~�l���ຼ"u�S9 �l	x��q����n�=t�}!�H��XO�0��J������x��O�}���[.9JP
��q�V�.�����$B�=�l��ƛ-�:|���`	K�4��Z����*7�#�6_&�`
yn�Z:�$z��`�lH.lN";)�_8#�qT���/L�N� �����T��gf��^�U��^i��6�	xN����k�<d{��u=�|5|V���9<`�i�o��:%8ͻ^�d�;���?�m;�q�疢( ���
��|J������o>�Z]_�����sf&!��MKm�o/������u*@~j���� �g�]�
�M�i�5l���E]��#D�n�ԹZ�kc�l3��S��Vsjğ�q�Z�
@}}Ѓ��>Z�'����=������
��I�hǝ�s��l�(���`�Ca�N"C�90J�R��Bo�)� T��:�O���p�cQ]I��0�Ȩ+�r��?�*=#Z��Eo��l��Z΄����I�w��ho������˼�/W)��N�"�\2Ӗ"�>`��Oߐ�Տ���u2�S���ٝ�k`8oeV��!���i��VG�q۬��HM$hm�B��@���0l���6������������C�G ��6��U�V��|E�Xn�.~,N�l��~傃��D�.�f����+\S}�-+�
�7�^�ML$��J�e�M�̺Ioҍ>�Wz4���:��Ē���	�q?x`hhE���~�(�;���E�^��p������b�6@����*PM���#���ݞx�9Y�Y-j$IxV�O�ͣ�P�/�G���
y��5��z+���z�>"��j��G�<<��;1�;
t�-qUP���z� ��U�FL?��5,q^B_�>:!�69��a��y5~�`������0�����9�]�&)�N�I��g�z��z�vY.�l�%X�?y\�o�
[��hN U!#���/�OD�G��*���7䚨[�t�ɕ����ɫ"�o(ۂ�/1>��`i��^ ��3�?��Tj:{Z�ߞx�Ż�m��0�ɵ�8��=$c��kש��)
0|��I�*��Ӕ�ǒ���c����TP�����S�w�@���
zU�:��e��b���6F�2}�h}19`�g�n�%٣�3��r|�>Bgvd�r�3H����_{�a��kLɓ���T��\�n���y��-�;��_�#�������ٓ��x�0�Y\� ��s>�u��P��oi`��ң@	���hAN�97c�	
v�(���� �@��_��lX�'@��
h�i5�M���$��%���^5$��χ玭s�۔ɰ,�?�?0��Z�j��2=����׮s�Bdb�f�y�o[�y!A�����!�g,�YF����c�tccS���
���H=0a�`T[�5��ڡ�
\.X0�г�A���QE��t~_ �k�c�&�m��^��E?D,��8k�}|#�o��
tk��i��i�`��8�i(瀹���L��m���UfG�2\0B9Ղ�}���8LD�_��v��� ���*�����ӕ�NLA����yoy���9s� �~���8/��
Wv5��=-f��������@�g���$j/h쭊�'�ױ��� ���8�O4�M�֔a���j��=�T�G�b
���M��z�ֶ.��bGɓ���xH��J���C��;�O\cÎ$Ȣ�{��D:nzL�����S�mc��r����bte�& ���-m1qH�'�u ��.E<�D��`gLxcxD��!�{�ABzz���#[�L�5��dB���5v�;�Z���A��4��ݶY;]�4�$*H�m�tح���^G�2NDQ�i�1��o���Ny���ǘ��E���@Ck�20@��]k $�9�	3���-E��d:<�f��-��׾�gc7oܟ�O�%�|b�ߘ�������5�922?;�������4O��� X�������fc	��$!YJ�)i�=je�%	TuӍΧa�؍-�Ƈ2�ިr����p�P��W�;.��d*kk�	"K���Y���@(_:e�xٮ�ҽN����`d~�>�<%vD�<,)rbtF��!���S7Er�;6!BR�E�ʡ�A�����Nm�`���k�c�~"��}_�;;�s���?�N�}�|%�f	(��5[+��af�(��&�f�Y�LX�TN=f���dnzh���\FTɈ�J	�w.�@�	ٔ����Ȓ3���}C�a�:�>�\��4\hs��(k�:�K2M(O�����0f:@sh83`�
R�A
d�����J�f��B�3�(R�kr��u����x&'ٙ��D�:�A���DN�!�������+���Q�v�A���> �¾�>�'3�F��'��S{��`t;b.�/�<Ye^;��h�Q�M��?�"y�PmE\8��-Z�2fYХ+�'%���oP�0 ĸ����a��D��m�+G=�3���)�Z@pս��9F�*�K���`4�XlxVHYEB    964e    1150�]���!��#~;b[��n�q�t!e�gZ~_���}�!��/�+�J%����^J�J}�&PHgDwVM�\?���jBm�w�q��o3O�m�Q]�&v�����]����i�D��!Ok���(����Qoj�k���,xٺWì'zk 7:v����v��h���zJx�����ē'+՘�x�X�O���?�@kn��Ϫ�+z��ѾCW���Q���!�G��@��p�2�� �3��i��t�H(�����r�f�����Cx�Ʋ���+�G(h}��l�� �HYe�s���"��P~��u>�9L�H3���ߍs�5��-���KT���:�=�N=$D a�6'�.��6���;#���P���\���bN8���%ȋ� �3F*^�	��ؚ�qRXeo� "���Z"l�d������ڨ?P��s��M��2��.��x��0�<}8�ǧ����FgB���KM�_���zt��˘�[l�^���4���`����{��&�W$�N�=������g�de䇓��l7�$��+(w;�V�!��q���Z@�?��}����T8�iN���7�^�&S��E�X,�a�p�m��S{�~�Wgɤ |�a�L
KD��R�od��>���R�Ĵ6=:�ۛB<jPJ��T�l�Y��qL���6�,{�+�ɭ3���8u$���t�͜�O���/��ֻ�6Yme�g�9s"A4oE���lA��1pa�Pf��k��lC���_Wp$��yY4/�sx"��v�&q�]�mWD�2pgI�m�cT���ceԕ
�E�Z��M/*	"�D���N���	| ���9�]A#��Z��L~������ 4�%�!z8��1�&	���\~hf�>|$���A?����a4H���2�ƻi* U��VY�?j �ꌀB���:�AS�w\��<�H��H�0��h��N���[$ZBޞ(���K&`�３?��#MA6�C����T��1*�f����`���s��X��E_D�iS�v����X��E�t,.��K��V�e߂�8Q�����'e)�A�]c��C��P����s����.h�C���Sx|�c�c�@m����y*��ǯ��.��J�Y��7���J�4�A��j�;�0�;?4�����T�����$\�C�*������?g�U�(�3��N,AK6���ˬI �C����$ù��W^������g�Baym�ʜT�:��V��w���8I�;1�Y�nT
<���QL�sq���J����abN�cO��*�R��o�\�+X���V:&'D��""�=%d�LP���uSJ Ы�Ą�
�c��Tt4����Q��4��DX���F�tl� �ԕ$�L�L��lf#����p��2<��=�)|�����xE�̝M�ٯ��LҔ����L��Ĩ��1N��Q1�)���OsX�-)拣���^�hv���	n1��4Kw~��URhr8��O�09$+5W���C[.1�M?�yP�f�w�Zn7\3-	�F3!B7v��#��	(�;7�g�4a��V�\�f�6�\��${�e��	�x8�a���MuAe���z�����Por'�fL������{J6dTt��j�s0�˱B�o�+����N��q�����<Q�n�av��gL�n����1I�Fpo3(
��I�?'������T1"B&eKë�*z�o�H�0��-;Pi�/�6
��Jʹ�F��s��tX�'�������(��ի.#&��P�ɑ�c��A�/���ǂ*��f�U��'9-��^���E�X>W�y�&:xp�\M��(K"k�C���JX@Н����!�@$p\6�T�V��uL:��\H
7��\t�X�į�ϨD/.�h�l���'�ȬH�����eJE~�f���/0K&t<�vd�#w��
Fk����Y[=�QJ�.Z�n�I�8`"��x��}�KvE�/��=�֢�	/�Z �Nm�m:�b��@
=��]?fr���JU��ZXU��!K�.��]�(G��l-x��1�	��TI�El�>Ѝ��z� ���Q���-џ0Q���!}�N�:�G�o�B>��l�Á���x�4�
�7��/i�^������c�F�2G@�):���6�_6̦�P��QJ�"-x���d��{L�8X�]_��
��iy.ck
mGR$l�'�Z��ã
�L- ��	�'�)�#o�_� ����j��b0���H|[�t��� 9^���������'��j�T5ٜ����S�kN�.���W�� Y`�p-�E���c�`�	�,�m9 �m�H6�������i��CD8�θ�kzO��� 6��`� �G�Y0g!{�*����;m8r���ѭ���;���������K���(&w��%��}�&v���^h�����m���-}��QV"��%�	z�щ��2U߁��Fu���j��Tf��NC��68xUr��;�p����%��En����톱�&a�` -α�����H�,i�%��ol��4�:��7��p���(.�{O�eN�N˖�j��D���s��W�^s��4A�d^���٥!�|���TD�ϧ)g��&ZA烃�&�����p�~��I�!
��!���@�dPt�n]��_*�� ^f�kA���s�mǹ'������+�����#T"i�`Z�L��A�s���=�r��o����[��Ԑ��i�pgJ6��f8q;�%���$�m���*���_��%������y��Q2��t��D��t�p��HG�jq��ia~s.D�_��i��aM�:#�j��Yv�{��_2B_%���!�@�A9S^� N�.�7H��$}�H�-��M�%�`�Yj�zw���o�[�@IeOޤY/�p	���k�#i�vq(ޯ�ҟ�[([��D��b�4��\!�B�JRw�&�a�(O^�Yv�E�-c��{v��ln�,8�gn�5Ji��brUAì:c
�~ZM�-���-U�ۑ�;�ghN�|协�)FZ]�J99�%�t���F*~�'6�j�0}3�p~�{��p
��&Iq��n���#�y2����b�� e,����3��U.g�T8�̨���#O	�"oV�F��A%k�Β�%x�V�)�X*0x�����$b�!����F��2�+Ѱ�=h�����*�B�A6� �0���Ŭ�]��Hu�l�'^EIQ��zr/ʛ�e>{�g���5�{�Wg�����B���)�7�T
�0ے�����q�Y�Gro51 0�|wL�$݉�똓p����zJr�
;�L���u.2�O�Z=Nfa1ET>��>�������U���q��N��m~\�@<D��iai��ڲ�==EM��3T/���M
��|��c&=j�+B1�
;��&`��l�����]���^���@;VY��dy�[ď���?#��8��`�\�%�ܡiխ�
lzPt�&9H˕g��b�h,�aQTR+�\E̀��n�6�x���8�Z&b�	�<Unex+İߢ�;��B�`��S+dJ)_W��7��Szց��k:��M��S%qEx#U�a��ye���_���g�O��إ�&֎7L�7~�H��ۭ���(��͠vU�,���6��f��@z+�1g�w�c��9	����5ͲVLmH���V����d��&�vz���<&G��tUe����JZq+�wf��|��P�L�D���e���L s:�簍a�]���C3y�G��I8�I^P	AO��x$k<�������| `qS�3�i�
���Y���^����OD�5��.����w6��m�X٧:�W�Q�]�4fT]JcD���.Y]C��5�v�g\�w���,&P����:��VeY"Z-'M*����5������-��J_��Յ��Hc�i�5�uL	�,t�.(ES��_`l �x�����u�l�c	c��U�ޒ]-��!�O���咽O������t:�G��#�πl���V�'�;c\�A¿���O,����n�^Q�X��Z �=��G�%��0�i��8yqW邆��կ�#Q�S��&����:)�Ty<�}B�I�/����g�ăH��B���{5���,���M�6���\�(l�`Iz�+cG� �:��Q�Vr�����~�̯G���R�	�.m�a��
�`�=Bcw� �Aצ�֫ѱr"��C�׷�O��"�%���t��8�3��$�ѻ0|�9p�V�o�p���j.Pp�y�5�qtdNq�.�C5��s��k�fA!Duhe���Z��R<[��Y��.�k	!Y*�sT��������<I
 ,�u#%9!�q�#��	�4	h�Оq�g踯t!�$S�ݷ�����#���3�o������