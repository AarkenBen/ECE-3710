XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���;A���3w~�>l{�R��F����g�~�c��Y�Y���,5K޶�Yc�2]iL�Kv���[�݇�U����nV�ǋ�q`_�ݚ�%��|�q8?��TMZ��Hº�OV0�0	*@�3Y��H����Be���q_R�Y�3��8�Fw}v�&�"F�x�\A�2�G�ly{��0%�O�� 7�$8|�^[Q8�4t�ڣ؆�-kI�����,h�~"���h���%�h>����~�%�l;���?n�����z�����S������?	8{��r�dBVJ�w(����xu��l���6vd�Ȥ��G)��_�9D
K��{r[�_e:f�X�#	��mtfO 0%��a�B�,4HVW��8#ҴGq�q��^뾀��-� r���Q�AK��0Y�ć�G;%p�a�D�'�l�_E�X�����n���sw�e��T��a'W�Wc����ؼ�cn����J�T��9����.>������Q��|a[�/��Fe\�Yy���&3��=��A·}�*�3��0����áQ�k��-�|s�t1�����}��u6w���4�a��������_�#��R�1����Ѥ�����U\����;8������c�2�a� ��hhf�,�A���@i�0J��W
�n���D�T��@cKI�؏��`ࢹ��Y�݋-�ښt;���/�>�w�N�Gg���$u�Γ��P���$�E@�׆!��'S��W��f�}n?��a�vv�=lA�,XlxVHYEB    fa00    2d60�Pv����K��Է'�I[5���dȭ.1�$&k�9bwi잾��ģ��a~9Jc �K�v[12*GZ�z�C|$D���,&!��<�^�
y�N󓠋Öۗ�6$�&Z�;������K��N+��k������`-�72;d
O;+�X���,�< �鴷ة9]ԥPv�J���Q�ɲ����,��ʸ���)##	��k��ىsV�$D�.lh��D��sW��k|@�xei���������e+{{�ӳPXR�������!O���9b"���8Dz|��>�f�wSz���^��9/��+��u#Ո;�"�}ig f�P�����%�uJ����]��B���.@�y��U���c׮p�g�!<������B�E��X�	�j̖K|v���-��Mn�tv���|���Y�_��~��c8�C)=(�eU&��"�(}f�$?	�lr��#�dw) �������!/{��1��JR�dIC��rDE�J��?�(��ې�����@�]
�o-�k#��pc8�Qh�������O�Q����rz�tyP'�у��asC��8f���������@,%�+a/�#���g>k��A��ʾ��s��e'd�>D]���&:������-+��
�xj:-`�*<<��O�ه^��!��7��lxH�bw�wI"�~D
ǽ�ꐐl����i�*������	L�ho�/������:C�~�����g������r�5�oQ=?����綽)'�����+�ɵ�c�IR�S�5�$��i>Qn
�x}V �� ���%��Ww��K���")K�J�tg��TB+������!�1jbD�B\�=�1�&�9;M�!��4x�����:1��H�w:0ƿ��\�F��R���c��~��M�=�CQK�A	}dy�=���œ�%�bT��
~��w#���lƑ�ˉd_�)��E}��+!K��j�U5
�9��B�U�5׺�[O��##�c廤��M|�;_��e�u��*�Q<"¤q�L;��M+w|r����;AeC:={�e��~�q�=nH�p��z-!��53�����;�����
�T(�W=�Z�#�������D���һ�.���L�P�	��'%��Z�����RO~܈���R�@}�5��1O��/U��Jazj@�G��E�����
��2�/���C֥K�nk��Y����Sk<_
Y(�2���|EǠ����,�?�X��8�ť]���R�+�B3�?q�{��J�l�R+���!��i�:qBɾ�Bo-�wk�.�JGy���+
7���R8"<����.w8sk�[I����'@2�^�o��86��t�)ם^��,ע80
�<^�3�����%o����+�YP��l�#�����$����,̊��$s%�S� ��I�c�)�#(������u4�T=M�3�v��*��ͫ�SL�LBI�_�h�5K�}�6+�b���19O� a!ý�v۝ڥ������z�ōC,W�}J��6�mQ�n�����g��Y���pD��|l�+y��z���6��ϵ'+�(�>To�u��@4�z}]�7�3
7��V�#�H��`}���m��I��B;�O��>���3Et�v�����4�ޠJ���dg�r�4F�k%���ZT�r2O��]<�I-b�F7gP0}Vp�${߫�B+V�W�Ӽ�5�έ׋F����@d
U���A�d\��H#A�-�Jci����v��>�f�B]�zj^���3���#A)(�?�l�Q�F22T
7�B�i���N 9u����*dA_d���c�?Y9��0O�jX\�mK�u������1R���nt�8�T|-jY3��ݳ��ˡ�����It��i<������4ӓ\�%�z�+ 6�ꮯVx���4@/�{���׎V�v�N�kg�w���v��]��Ùo͌� �Y:~A���EU��':��QU���ʹ~����۱ȥ�p��R2�E�(+@�T�ƾ|o���W��7��C��P;PG��K={tl0\�זv�8��u%:ǶǠ Ч}Y�t~jq�ê����n�ˈO/��W�b��r<Jr����p�'����t"� ?��?�7��h���u�!������ �~��lQ�s�b$�<|=$�t�0?!9���C�xj�Q$v��1�G��[�*v�MRi���\���&���n�k&�؍� �r��e�,|������!�k>�C���#�Q�X+��0=6�;�u5��~l��>��Ku�z�и�s�����g�H��܁?�������������U���9«1�ڇՏ���<��)���~�Sv�T��Q��Ip���	?�(���,��ߚlM��x���P�h��M�+��u�
]2~�?�;[�(w0B�B���W!8)q�O��"��F��Zar1���/��.�4Q'>�����ω�1������@H��P��������iP0�7����y,B�_|A�C�<��K����oP��'<�k2�i�3S�&��y=�	^1��`���7�j����̘ID��`�O� �)f<)���c��BĽu��P��.Y���R�<o�<d�v	&����x�}�N��e?F����X�a�i�@��~���*��>K��� _P0�L;/�u��������w��Ñ*/v#��s�n$�Z��s�u`Tw7z�B�W� ��5����O���c�M"�%i���s]i��3a�)(����z��qn����w���rM7G�
2_�+I���Aj�0ˤ;�����n��F���#b���Ÿ�T�\����v�^W���v�}�{�m�ޖ�>%1��;lf��w�o��$ۦ6QL����݇'	�nO��5�ܐs����dS���)��`����{ oz���� 9�7J��mV2�N;S����P�9,#�TR�|`$�"݆D�˝0�1^��}��^W��f����oa ��:-��M�����cy=T���w�}|��*̇�0B�ys�}�\4�ߘ�#���M��vr�n�*�y�}���:h�7\H��ԟ�X�]��/Q\�ci��l��U}Ʋ��Q����$Q(}�0����2a��N�,�I_b=�"����ɒ�����H\�U���nL�-���u;�fй@���|�Ib6	����j�q���,6�
�ݝǶM��,sѡ�f�9��n%�jGsiLD��@3&�/���?�\/��9�I/��|X��7�=��}4�0	u�E�ƫ2�\�5�n��U�yȎNJ��Ԏ��*{j����H{&�3� sU� %:$͕�K�W�!�AU7 ���?�+R��#R��|ʆ�k{�B���{I�Hi[ v�e�D�~5 U�d������a
0�%jf��k����X�OX�m�ǽu�=,?�0ffa�ۯ�k���G�R��/�j;�0����9k?���7f�'$�q�JciN ���W�� &H����<�>;�xjYƳQ����JMp^�7 D�p��-|dt���)E{��f��r�.�nLA��L�\�OwG�7��Ԃ]�[G뙣�� ��8��U9Bg����mV8
�fSL�A�J%���oE�n��vv���pI脸 K"��!�;3�J�+�K!%c�;�~�:�BGHp�Uzs-d�J�UR(�j�NzK#a�m�Z����Q�I���l5�w@��J�Bt�1��e��HqsǗ�@3�r�~ �c�5������q?+}&/���{i��6�K���O������tV҉>�yXx�\h�j��~�(�f���7�f�G���8E�.m���H�Kh5���S������3��,꺋��>����i&��0R�r �˸Z�+����A��W�@��+G�9w���յH?��<���-����HO��Q!���(���몷�D{f�§�=z��;7d�sج���1V,��v|���9�*h�v�7Ct��Ȩ�����TH�Rџ�3���x�?����a^��^��w��FyA\�F�h�e5��W�5b���M���w  �_'��ߚ�6�o�?�d�7��&ǐW��P�A�s�j.]�b�B9�f��]B����ێ�������H����D-{�}ph]~��C����'�B��H�dnoj6>l�=�P��l|�� _��R���Y؍Btf�_��o�(`��]Ls�|�(8��q���8Z�H�Y�4����ї�T~ S����9��uu3O�l"������Ǚ��vM KqV8��|��[e��J��+%(�d���	�3��i«��.�o M�Զ:�f ��V4���{��1��J�d��c�������X�U���Ie�PJ�7�O׳��lFt�D9���B���w8��$�3�W��T����5 ����ݤϗ�$�5/,|�]&9��L
�o�/�>}���jU{:$��g�X1���q�	���LG����PVsN�Gv��cwo[V:=X������]۵0�Y��1[k�������O]e�M��\����p'��<�B%J۝X��!SS�T��~�pp�t��Ō�����~���|�ٞ��躤(ڨ�G��C�uV��ԭ�?a$�3_�B���s �;S����F2e�����0H8�SU�$��$v��&��$�6�
^a�BrDmeG�� �_�س�n"���ζ��-�s�bj��I�־�l!?|#2�m��eϽq�:h#�(5�<���b���fD�B'��8�� ��{��r���c���<������	������߮��TᏨ�\.��K�v�Q��Q	x�v�3̛��C�IN�{���g[�^a�!x���������:�ॐ�����=���BS7�$a��8�#�؁l���&���ȼf���S�M���@�T���u�!��u��0\L�*i���H��ض��h5�e��3��R��-:A�R��R��	!���	�>���Z#V�LW�Pn�%�&�������j�,HK�;�C���'�WF~���`Xv�beE��o��JqM���
<O�(�n�f_���?���>����AK��; �5� �Bt�(� �n�C�ʆ+&�8�D���J	�M�$���q��"hr�Ei\��2���Ӡ�pI���D��f�{0���Z0�,9����:dw'��/@U�DBE(KИ98%ņ�-�{"���@����Y�ʥ��DA�|����\�G�C%��+}?��=/%�z���I�i2򕏯�P�U�@��2�|D�<�"x���W�L�V����P✠q�l�]�N�=Ђ�r�y�4�,�S�qԮ���)����%GO�)�/���JY��q��D�k�s����	���
���(��c`��T�(���,�N)*�u2r�ײ9�%���k��0�W��^��[V�R`�Y~���e�5%��:U���`f�.��޴jϐ'� ��ar�R g·�P����E����ry����9�eCc��8=w��� ^0�]�`�h3�G;��$j��PH��`��D�$�h�t�M�a�3	�B�Ļ.���^�<Iz�λi8q��
_�T��v�S)ʰ>.�&k,���K������9��S-���Wf.�����W�(蔞�$��Q�!Yf�ѫ�%@�M����`"�:����Dyk�pG�#?��p'���K6Đ�뗡��#nph9T؉�(�
�fk�U`c�S�ē�������-� }~dT�C� ]��2���C,��1ԥj�^l��䪼&��P�C�����H����W��K��w v���0.�	���?�Lj�^��nU�g�.���lI�����]���&������&�r�0c,�����K����-=�r�v���3>���U���?�s�Tu[
a�Y����2q�n-l�K��d��w |����PHA�c���UL=��9�!齝HIa�s=�)H�<f4,]��
��v7��e��XJ�O<����e�S�;�ɱ�����w��4�KD"DǷ�z֋�,��t��\�}���[?5K�/��hyy��d�!U��H��[�ǚ�^��b��2W��)F�K�.�@���U>�L�j)��&MwgǓԑ��w&�)YɤP�ǂ�R���b!~����Uᅟ"������^�0)���4����`5?�],?��祘�ڳ��>0=����oQ��oK����C����s�\��}�:�+�ݼTH��j~�I�3��.��&�i����ޑ
	[dZ��{�bqo0��?�Pd���Ir��^��E9x��Q�s�o�?m���9����}~�J�P�רzf�F���୐E�����'b�6Ӊ��DwwI��$fU_�����[�t�������= �-���
Gk�t��/��y7ء{�$�?R㲡��*3�3bpTUw烌���"	��O�����	$�xyH�ɐ]��q��e?�	� 71�͚��3&�=���8���HF������,$�	z`u[:�D�8wؑi��v[R֤�'D�����@Y�h���}�
)r��y��M���z%.��3�SKcE�Ъ�y�����&%�$nC����k�>]%�x ������SGj�[R^���c3�*]L1����
8(�؅����<k4!H��^a=81ؾ��P���<~i9oLY����."9v0;c�<ͦƂ�����7��pb�p�>(gN���e��l����[7C��y�KZX����:&͖�]3���Ou3 �1�7cR:����Stű��XKvG���^#�"��
W�$�mY����_eu;�t_>)pw��ʻ��h}�p���7C	oa0���Z-�DD��2i6��P��U\UK�4D�$���fT'��Þ��f`���.��t�C5o�3��i�Z��:�A�l�J(���Q���pyev��a���Q��ۆy��Մ���������������V��14yq�A~j� :N9,D�v��c��:������B�9�e�ƌ4�!��ZG���<(7��	���4I��:B��2)M���3���J:C�dذ-/�b���|����/)��p��~�i/ �,��J �[����(Me��1?�x_3�en���Z���z	�,�e�@uSy]��<�9/�&�OH��^)ZF����%tR�0�����vES�Q�.�ڐq%Ԩ�3��a�q�
�z��p��!��������mc�5	�^�M�-,�Ny%T�"�"̌%�p����J$6$�b�]��g��bD���z��墜�L�A Tz�O�.
��l�`Nk�d̆+�c��m�+��7N�.ٓg��5��g��>���P:��*d�Yc��0C�c@��W�e��{�|�S-s���|��}���Ȟ2���P�ݬq�MT�d�������gp�*ޝ�/���1�:5���1d!t��o�n��͓�[�Q�02Lȳ��{���ư�T�|��q���ߓ]�%v�[*@6A����3��I���A�W���!n^������I��.�oU\Z���Rxfi�ږ��|����j�&hN����I������,�R�f���>u��G���6,���ȁ���=��)|�G���xBK_�o�����&PKAe[
�E1a�B���%�|��Y������7��N2�eO�<����f<4��P���S��n�m?pco�{|�s�����ZXǤy(���L@��GG�I\tY������!ArV�ȳ���M��G�Ze_������;��4l'
�Sl6S�
���g�����v��/w��ڲO���L�l�0$@����_��S�p����M�#=Z@.%PB{��鞏��
���~[z�r�ռO�`}U�%�	~����ŲZ����JhILMT�` �$�� qF�ஸwE@�$w���B߽d4F��l��*)nzD�2	'���˘zݍ*���+�H� y� ����X�����h�����S��;� ��_$gF�%J�i��z�I��S�Ԧ�1��O����'�W/<�n4�@�Yze���2���xS*c��K����B����}�K�k���\�,��{��?I�S$��}I� ��8|4Ĥ�����mytI&ZD��pAjY��%�.��s!C���8r3Fyw�<�{i�Ϊ�f=3�[�2��y�Mօ�����y���Q��~8����0]Pϭ�SPR��o�����^CȾ��{ه~B(P�9��)O�N�$���ҍ�娐��	\E@����G�aŻ����xL���C����V�N�fmmz
V���c�BA�q�)�r.�:Vt��;���0��7§�u���st�vH��@�D(+X{�ĆOP�j�3�1
-�~�W�#{��!ĿO�2M��k��)��)2��:����֎����Aꄴ�ER�<��ҟ�]�m�Nz�Wj&���N"Ň�K�W�ńs���q��[d�u�;e�U��2���o89;w\i�����#U�J�2f%V�ݤ�i���?x	G����.G:�#�)(���?�EZ�lc���`���Ьr��>�7w�O.?5��7�!��喆?KrDQ�3Wڇ���P���$�Qp'u�}:4X����A(U����2ʦӴ��ޭ�,3�X�-_�\�I��?!��$���M�e�]�u.	��u�/ɝoB�%IԂ��>�}�t��Eo5I�n�Ank��6�����v���k7Ӌq�C%Xq�6�'��@����܍�8�������|���R��P{F�4�j#,�&{�!m������w�3b��Egl�%��O�.c�¹���������M�)��Ia����&\�0�yd$����G���=��j�9�u4P3�fe�)��z�JߛR6i~���1a��Û�)׼=��#Xؔ^�R�Joi�G�'����^j:+�9����������o���dw��0vۋ�"VϢ��X(W�/��	(q�>>��ظ��s��5F�������,M/�"h��Y�Q�J�AHTڹ����E��$��'��nl�V�?O��=э�'�[O�K����:BBy�sP���H�:l�"���[�#t�3�ᮞV��������,@��ՙ�D�u�#+��UZ4��pS�&f~�@D��1��r�a�!ad;��Hn�h
��1�c�qu���q�b}c�`�=*�.X�J�";��d���� :���%Q$T��@0"L����Z������c���6:&�AޢqJ�����<����j�S���1���&ul��z�G�!:Ԡ��c�$��3�]�bJ;o��S�Α'�KMx���b�����w�J����9)Fzx�q�0]ܑFAX2ԫC�#�R�A�5��e�i���I`Cn�΁!6<��c7!�,[2�3�Nlö8������=1&���ۜY�\b��8��mgD�{l�o�'�nB�!�T���H�";��� �P�{�[4+��!F�r��x�5��{Jb��R���1�~ܫX�Z���y�B��V����e"4������gϩW����HM
?�e���%	�W�j��E>&��馟*��b&L��ZĔ�f����|�o��au�6@��ز�^ĩ9�	r���U�N���N�̎��	:G�Q�P��+֭I��訜8��8ٟ�<J�\8��_Y��R���J�� u:��8x��]H��AoB��5��g	��`�@�@��-s�㍹�i���߿J�~�y\oh��Q7��3�*�R��@���@LKi���S���VֵFȳ�4;��� ��ڸ��ϋ����]���tQ���Z�ͨ�wB1�?�����$Uu�':�&�,Ii����e|�v�%~%�A���Whc�"���%5 ��_��[-�k������Os�g��3��DY�j�yU����5S��P��L�����}DV�z����2}E������-���BZ�Y� w�е���?�~��yVI�zJ��\�1ص։-G�0��<L}x�O�2�9�GS�7*�@M-��U&���6U�%�N�颃��+�Χ��1��|�P���xua!k"m��Ԁ�1�YҮ���e�SOK"R�r:��5< �>�s!��+�V�s��-�~�nS�x�߅[z9w=����]�s�d��G�tH[�Od�9y45�Bּm� gm����8���M���ғ:6�xX���~U�U����䩂����iGn#i�u���{�&l�>�9i�7��\;J#,�z7mo�vG�y�^n�:���^#�͍|�B���8�r֕�����J���+��n�t@�xཋ����[��ӑ��P^������d/J|L��v:��N��޷uQEJ<�4��/zc�yT�%{aH����pt����B��h�-���"*��"��k��ΐ��^Aع] �	C��ć/{�;驪{*� �����͚f��\�4��+Q����	������ȩ�L7���lz�Z��%A���*92g�H�r�(@e%d�-_��:�z����f0Y���`�#��0\ύDxhG�d�ˌ�>>�b�g-����X��v~�"��t,�}�Vۦ�'D;��:����A����dذ�#J�� ���l�c\�gT����G�2y��g%כG�1+�"�n(��8���`+���LI��d�ЭZ�y���X[
8�8f�m��6E�~���c�%���m�C�z*~y�j ��$�R�z��M#�=�N��~�b�6�϶���"򝵯]q/��p+�S���[�lo���5)rK�Cnr���p:��j��jl>��P_i-Рo� ��f�8�EA]��u+gk��D���:���B/������X��Y�x��(>�x�@_PJ+��z�0�'�AK�e�b��m�ND1-d�q�B��M�'?��u���>���^N��+�P���yb��eܚ�Ы��\p$���ge!ɗ�<����|�/��*�-یb��F�E]�\f%@�D��-A)x�����_�F����:�±�N�}-���������j��7љC�$%�%��(�%���Q1�?N�����Z�~ٮ1������J(����s�t��/�[��5m���&� �δ�yΙRK���K�X��@�l!	᭔���O7y�UYY���c������L�&E����3YlA�ʳ)���ߨ{��`�Qr��{$��h�Obxa����E��~t��ᷛ{j��y�/����I������)���>�Up�4Y�IH���C��onv]Ԍ�3��S\�h�:��c{��� ��Z���9�R��O��u�6{��P��|�S�{�U,�����N�d|��3f�<G,�?����HG�h�8�y�R�P>(�@��'1�ι��n����(�0�F-�Oh�Uqb��V�Չ��)T��R �,�o�_�|+�jBt��"��DrH�|%�Vc4
�B�eӘ4��& ���vJ�j懕XlxVHYEB    5914     f20�|����T���ϔi16_!�w������4�􉜇M�Ȏ�;��X�<.+)F6���+�Eў6 }љ)Ʊ�w�Mf���XlmB��a���˹4&���Ln�w��*^~�ѩ[f5���ac!Ϙ/ 
ܲK	�,����3���NG*3h�B��p�̸T�`ϋ	����cq|X��|P��T�#��@��A�Y� X|{E�?qp����I\g�����Ǘf�WE\�k8�7���	��������� #�x�s ]�y����b�D���XgG�3VQ�m9�pD�D�Dǅ�>�������*��L1����a�2���>��mu� ���!���~�(���|M��(VY��p^TD'�� �E��Iݖ��ݍ|�Kd�0Us�i}[�3Tů�ߑ�J@���b�9=�gi�CfU��v�WM�֒rU�}}㙎��GM�[��Z��M~`�d��+�ܷ�"��03$�w
�i���yBQ���a^���o�B.<
d^��� �E���w����b�Րi��~�ei���e�y|ԯ�
k��DO��Z��R݀�[����U�1͕��Y�c����#҈�"HYn�7�IwV��T_F\ը���d�^Me�rt�L�����Hހ?F%����!��H�P�K�������������N��+y	m�V0<�;�������vG���O�&k\[����޻�=V������M���Q,f�=��8�nSS�Y&4ȋ���qQ��
��ў�,���ֶ��UI�@���{1 Ư�9!� �rU�`'D�F/���񚪄���K,A�:�*��k~#�b1A,ŗ����FS,n+B��{P�a����|�渵HO#ة��̇n�l˽�ձ�n�i�424�Ų�W����5�}D�~,R�U�r��T�V�>M��X���P�!���%��")���_ˑ%���$�P,��Nl*�B{�,��y�]%�U"ߩ��S`Q��0��^2��"|~��@�ǔ�Z������3�<��'�-��a��|���������9��9E\��+�y~Æ��+
�	w�52���Y�aZ�)��̊Rk�;e���I��`?��˩��� ���n���Z"��
��	C�n�{?��$�|�����D������P@��ZFT��@[l^!n��vi;\*���Wg��d�k3<W��y�.]p+��.25v����ey濁��AW�hP)Jy��:��X՚厈3Bj]�r-�͓25���"�S:�rx\�(���l$�Q0�f��*T�����b�kl=�޶G k|��۷FĲ��ct8����:����y��E�L�,�-Q/����j��N��[��Y��̮5o-��^TN.����Τ�5�C�m�Rʍ-~Y��|��0R��h?�$��L���r���j��
�[��c��Ax�Ϳ�:T���۟ڃýu����
��1�൑0���hofw���hy�lP���x#�鸳4~&��$m˪�Mp���0���j��%t��(����iwf�|/�4��2y28~�+	�B3��������ٗ�S'�����T��]D�R��	Xv�Y��e-y�c#i�R�����ӲIL�N�\4cvh'6�|3nI^��Y^��t��ZҨ�rR�D�	�lt��1��,�٘ݓM9����'jU0�i�u~_��.�����+�s�6�&>�h�J��A����3������>`���eL�
�#�����ɶ��ьZQ��?V���Po6�x�j��E��=�(�Ag�(����E�2o��X&�L�
��Xѐ�fz�����J��-�θ� u��	��,$ǲ7r<.���h�.��v�m%XE=t&���}s��O4����F�ny���ޫ����߻������Y�=L57������6ʮ `_�c^i�����/n�OIu'��w�@������C�'����r��I�����И��)���?%6���V]��T�
���|gS묟�Xr�-��P��$������T�Co��*
\ �͜ש��-����[�r ��Y 0�z.@^��?2�(�r�Z$�6�Ě��4�~��c��&��<���Sܖ�C��d���2�er�QTd�d5��8�4�&��6����l����Bw�3
�q�Bc+�&V����Z�vkp�fj�29���;j��PW�ۢZS�a^�1K�������v#"ܞh2f���F>�D��)�Z
��� 1��6��F��V1�T�1E��3�����J	G�KW8��qѶ�'���8`�mn�I���΂�t�=|v(�R�\��GU={���	LJ@OO��a#��2�l�rJ^�?&��8��؀��&��S�GE���Ez�j��o��M"�d�nI
Q%�����<��� �ֹ�Ec+�o,�%n�����oaK^f� ɟ�\}�e�\#���=�Ը ݬ�0/�+�=��!���%��j.2��L�dG�P�ή ̫G����,��O��^T����j���̣��u��9g�M���Ja�G-�B�]��]� �74h~��f�v�qU����C���C�k�g���'��r����znG`u��D��`��(6�����^�U���#�|�Z(������ITz������x�p(e��K�|+��R�ۅ>s��?�1m����2�A��G��d��+��<�-ݿ�h�;�7	�-]��R�XЙ�oE̓ ��i��7Cr�cQ��+k陟���=	A6DB����;*F_�� �9!�ٶZ(<�lj�rTb�e!�a'WF�AU��è����2t��|<
�������T��D;�!��|�4��'������qj�=�=�q���yrU����qAL���9z�W��>�>��{��i��3��,�c����9Q �lԤ��v�a�!T����+�F�z���)Ή+���b�`iOힳ��������T�F~��i>`ơ:��7��i���z��}	�����nMd�ȿ��J).�*����f�J��@x�Ҧ�(,��3���- �m`�����toVpTҾ�����TLS�9�)SL8��Ӛ��{�DZ��� ��ms�idh����/"��=;��i�@f�lNj�ä.{[������2��e���+�=���6�t�}綅�������ZJ��<܏�辟
�!I��-�m��;�O�qZ�j�W��%��J2]�w��D�9�$1a��a����,��V~A{�o��.v���Āҝ�����L���kɽ�����bSgz���NcxE9��|
������+܈;� �����TP��U@���R�Y�h�M�
;����� [��	�cٝz{��	I��75�&�����gH��C�+ ��%Qq}���o�x#a��J5z\Р$��� �M<��~�R����\�Vh>�P/(�� ė0� qEx���%@j�P�Zh&t���+����i�\���b�u����{p{�A��cM��j!Խ����� �,��͌g�����1%��#r�W-�Z���[�b��������߈��t�7N���O�q�6����[��*�q������^�����a�X4�-��3��f�"ۃFʆI�,���F��h�s��$���]7�$�\��{#���ї򵈢,ى$|���ɣ:�$/u��I&���C��loyGࢫ����xf4�c1��a��ؑ�2:���j;�]Arw�;(Ϭ��'�:^�tq�H���y��_u]3�<C3hF(7j��=�Z�@�