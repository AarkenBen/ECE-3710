XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���^@�P5�I�C�B9��S���Y���]����CR۰׽�W��I��dHJ��~L{�ߛ�/��۰�h��+Eק����.ɣH��O��|��`@�7��@�B��/��_H+�&vY{�_ķo3���ʊ⬽�o5�:�K1�I�)!N	B��I�g�0e�R2LL��a9������܀��p�/�盇G��)�bП�!���3a�&1��^�xmC�F��v ƛ(�V��0~uu��ڟS+�Qe�N�o�l
��a�ĺ�َ���?^5	� ���-�όAzOH/�M���z�	\��}�*$E}.iQY	��V�KlG�/��l�]�͹��%��G�b�g執��v��c�,s"@Vg��U����X��^E����99XT�8�;7����z� �[��֢�� �r0�Œ�����Z��sLO�,������|���a�ܸJ��FU@�q��dm>`����1ޜW`��ۜ�=H�.�bpI]������)w�����4Z��W �?��Ai�. J�[]����s;*�Ս,*v���K)�����4���>�Fw3C�������*`v,�.s��&Cޭ��D$� ���#��e�H�m�c�����T��~44�����\�?_���Q�E_E҂��$H�;u�|g�\�R���C���"V;���.�;�#G�P�A�S[n�f�L8�Mr듬`B��&�u�jIό�V�
f�;��*�H&��@�í��DIk^�xt��¼�V}c6������G�ڕV�,H��XlxVHYEB    fa00    1fd0�hF�~�������;�������a33\7�b�U�+=�{�e~#S1gˠ;�R�-,�"�9��oNP�̾i�P��
���y ˇr���_o[�ܕ�6u�yLh�6!��)��w�a��Y8�[��!�YsNE&��l�ĝ��ӗ̰2_a�5��I\�3狮� 5�a��~6�u�>l��Z�E�����z��a�B/�D��&֙��c,z�t�M�l��Ɂ�0ZɌ�8��9*����!ۈ�B:�V�z3O���A����Ȕ8��ָƳ�K��T �:C"����]�(�/�M�����U�����F����s*�^��)6��7ŜZO�����&����h��Z����2�D�.�m��w�:>��|4��'��gΌ^��Uͷ�5��|���o٦<@`��0��7۱Q3�=�w�Ѫ���)-��J�(^�H_�x�����<�($�}#�	s��L��_��i��_����W"���5�ׂ��i����}!k�/���Z[=��KW�ф���	 V��Һ�B�]V����	�1��_��|bQX/���*���� �ǒ���za܈��Y�.X>��.u�ː��Q0�j��d�ڽp�Pr���^�"���vYlw\Mߠ�o��I�G԰��%��o@ή������E��:ȍv�V����=�]`澃!1��ߊ�=u�bO�bRr���B���bi�Rlx S}����gɃ"���RL���ќ��atpLk��0`�TL�f 
+��J��kHe���®¯?�K�;��iOk��тΦ]����>		�z��d�|E�C����ɲd� �S@1}N�9%�=�8A��YڝHkԐ̓1j}��Ms��R��2X�������tP��7g�,d�p*HX8Bo;}	%�O'v�}IHCMų<����P���([��Q#}��-�y��u��"bD�S��7�Qj�D>+��c�T
��e�\̓�+��nJI��'��	c:�0����*���@~u$�S&@)�����r�^�K�I�r8=lLᤦ>��{n&����˗	��Ju<H�<](�DN,�>[��j��֖��S�Gu2ԤFSj.ko.X�+-kZcV�h;�iY�,
!|XO�=��!�����={X�k���D#I����y��A�?�l����]dv�k����IgD��A:����1]S�(:d�K.�zr�/P. ڠ_�B�p�m{�T_�7-2v9�qM���n3]���Rr^&�~�{<���Ãh�n��	�B@V<�������#֋,B�#���Z;i�XX���0��2d�=����6~�5�����_#�|YLI@�A؈4��Y�&1�ʮ3Y�����/6��GY��/�	h[��L5n��6Oq� ꥧpE�g� ������E���Ȥ~g}wA?���W�_7M�2����aF'Fq��G�* &�����M�~tt�8��{{KY=�F=�%���Ɯk�O��t�t$W���7&�D������W��@צ�E\K�LՎ2���"5R"6*o���U'p�O}��E�.Y%%y��a�-]��f���G��eI]0G�Y�KY�i]>C�PD$^Ku���C�B�W'����}�E)f�z��������+.�L��o1:�Yϑa�-*`E`O<m�qZ�Di`-������Z&�˒w�K��c�����:%Ƙ�+���*X���E/Q/)!>1�ۮ��1��=��XR�xT�����j\�ճ����KKb����x^����q�t��rZ��Am��[+����a�-o��<n��L��(Cá����ĢG�!/?�p��	hY�Zk=r����2�%%EU�T�h��G��ML�oi|C�?K�o��@�	�)f�:` ��R���\w�2�:H� ~�"EM��o��'n�W�`�����M��|�Q�_�,�8�&#c7�s��/��8!-�L|� ��L{�P/���,�h��q�7@���V��U�Ԓ��qd�{l�?%A(?ɭ�
�"d��3zHU���,
�����@O�G]�p�?��D.�ˍXRȹ�ju��Q���Uަ;y�����)8\���W5ߖ��q0�sM!����ޫC�h�Z��E#���Ɲ陲�� �v՘6I�o�(�1��tٺP_r� e׀�����S��A�ơ��5�T�:Q�4�r��}��Ex
�&���F&s��2��� �j�8x矘[�����۽+��S�O	�ь���5 �Wԣ�с��~]��2KR�\��D(e��K=�?����@\T�s[�5S-�x䘚�9�]=7�i�Et�_�����#�o�r���b��Pۥح�� �|�$*j�������o$,�҈�zR8������B��平��6u%*�i���Cjr��hթIV�#�#���*Q�MgH�Z�#�y$�������������L*�g��C�CFץ�F��~FT��𯹼<gh�A-5LJ |��`�q<�!�k�����A��O%���T:�t�7�$�~����e�)$�M�5��+]5�o�Yb�{\�H�SF�'�����-�F���N&!)a3�M=sv�I��5[E�\Y��Om�á���?L�6n]}7�!!��_
�
�]%3+�>���r*EB��+���������]�i��>\q��� j�r(��Lw:X��W����a�-��#W����?��)\�;�'4 �9:<��J�wU3��yƇ$��G��Zc5 �ip �q�f=&ҍFv���������3���&Up]�����W�x�
%����M�L�D��m����9���^E���&�kX�ԙ\��$��-փJ�4��"�%���W���X~w~�&��#�ۜ#�ޭY���^t��I��1&\���F t�h�������TmL},ђ��_x]���UBҿ4���7�򯛘�tK�����t���᱌�2�(u�6�j���\���G��K��u�뱽0Z[�¤�d&��[�(�~/~(Q̟nq���/�x��4W]\�=Pw�8V��)�W"�עi�AS	�w42�yV���$h�2�̅(������l�g��?\ޒn����*���q� ����HǪKL(�
^rܞz9�e1ɋ���nU�J����������Ƥ]�_�1�ސ�����>�!N�m1���]��0t��|P����W�<�Ǫ��$���.�x�W��jζJ�D��)�ܜ�e�"u��Q�Uơ.W�Yhc�b��g�4=(�6|��>��ɀt�����g��Y%�Z�ѡ�����A���BF�ι?E�����*�������"��jx{��x�:�!f���V���j�5���L�7�8�fy�,B�E,�ޫҰ,���]g��BV�Kk��ib�e�+c1	r�US��7��l\f���MdY�+ўn�z�:aH�H�P�/[j��\kM7�x�,�>�!��EJVp��C`�@��� ��<�����0uhi�������{Z¨�'�യ��n�}�LU���Gȋ�j3l��V�X����p0hs����\���dvgmzb��s9 QV=�Q8�z��*_"�3s*!*�d�{��P�֗:1���x��mg��2"T~r��<{`60�ݟ�g�K?�y��&f��%b�k��\�K���#���Ӵ�xCY�1���9����q���rw�}�1g��=:d�du�!�1p9󖁤I4h�%q�Tb /4�j~�Zw$0I���1��]�Ry���B�J�������7�y�@E<��\�gT@[Ͷ_�ݍ����*���3���@I�:�����&��	�}�x�q�%zЕ�酊cr/21�y��#��SH��YE���vE�4��<�훴�s`��D�muG��$�,~���}��z 2�����Ax��N
�hO8��i���2{�b[N�:��V��a����`�cU��.���&5M�>'j e�#�T�����8�e}����Q� R�
s�����N�yI��A)�QկWp͘<)+����|����B4�?��2 &"[���6�@��^4�b�9Pg|�����Jy#���B�m����j�bD��Nj�W,� z���b�.�Tq
�aLbN"�]�.
~����.e�{+ǫ�
��0����#�Q�'-�������T�K�� �(�[����(#��۷pq��h�g�e��*�g�,4~O�m��0�H���_��ܧ-�_l| �Cu��P�I���j���SJZ�*&��EqFܝIsO�����" TAQHe��ߥ��͂K�u�LnyJ�����~��q���ekT��E���:}.6#zi��&��~B�0��K_%�F�����m[gTq�B&��M/��&ǜӁ��~Cgl��-�6U��m$SM����.�h���R3���.��,��*���X�V�(:mҧ"���;j�oV�k�0q��SG��p����(eO�8�!����ݽz��
��n�9U�:��\a.>m"��~��B�m��`��ݡ� 9�5�W-/����Ǵ��bfCF��@���Fț�&�k����HB���s^��ا���J���Y3ת��җzr|ε���俗��I��l�F�M�-0��aNU�3��TC��ч�_��9/�7��~L7�����-w�4$�8��{W3QC	�)��|NS4"N���U�o�����{���x���z�iN��)̓]���-��f��G\�Ѧ]���"�Gd����u�9E;���u<���XBW�R�<4�a��'��[�e����q��Q0�gϚ�I���"eHn��|y�8nX0�����g��H�+���2P"���|x!z����z>oʤ!�ײ�6/�*f!��Ҽ|x4i^*��Q��, �K��#�6�:�/ʲo�|J� '�C� �/k����+@�E�	�f=��i��uC�&�%״vi�)+�� ONuӡ��"��*_EH�p�/v1����b��|�Xgo����$"�V V��f�R��c�%|㑍��_���kp�Mt�Vm���E�9��}���|7��(�7ԥ��i�����.����~�����ײD�����v|�$mlE?$�L��|��^�r�r ̓�c���6.��c=�+2�q\*A�߳)8��y�iʻ#���(G7Ui���D%��%C��V��R̽���[w�^�Ai�Y�H�m֢#$�I�M����d����ei�1I(#W�����rTlg��x*l��4\���]����+E>�>�`$�AeV<��ʍǋ![�`��	F~ym)�o���/�+��n�6A�;�dh9h�GE�w3L=��{�me�i�F�G��h	�;�̷��0��l�=s��Yj� K]���y��[r�"~�,\m�ك�6B+�������h	�)����fn��h���D-��T(��)�e��N�|�a��+̕�l��X	�ƴ��^I҆,��1��Ť�A���t3�_���-Ey�~��EY�N�p(S�+����1D���E��ӐǦ�8i�Ӵ#s�Mw-��C��f� ^�`v* �E�Wz��5*��0I��A��D��(��Y��յK�g��qLG��<G��uz�G(Puy�Jq=�fO����3���G	x��B����_�n��r�M��I-�7\ވ��O��-�����l�̽�][�]�iG4����iJ"��$#=� X�gA�r�7f���6��3�W�b�f%������R��Ǳ=�[�#b�*L����*�S�Tֿ�,�)�[��,UT�c�����!x�*�s$ܑ�'z�KMh0�n,T��/��B�8����O� �<F�l�>�,]�__B++�9��q��|kF<�/�Zg����D�7�f��Cj���g�)���{��uŮ:��-검Yc�X�,�I�l8����-(*��n^��*rD��,B�N|��:x/ْ2�1�%ȓ���I���R%��"�[�c��x��Z.o�����ʴ�����iHQ�
�S f�mV�t���� x�?_���$�I¥��R�����>b��=>A��+u���h�9n_�����(a"|���f���z��I�����ѫ��ܮl"t��[);�Z� �&-�<t��MU*h��C���͂�l ��7�{Gpb%� L`A��KD�n)�����Pָc���>BAJK}3��òK}d9z�|?�g����Y�!T/�������.tȐ�u�'��I�e�g�#��޳��'[	�n��S@(��L�U!Ԥ@�o�+z�@��	!{W�9�2<���D�ت�����N�6��i>\Vr�A�o��f//�Pbn�\��e�/��}��T�K���%ƴ~�,r�7U]�T�J����ձ�)(���-��u�����S��JiB���A9����g&_�j$	��W�v�����c��u��j�E���)��Ы�wڪN��|H�y,qQ��
�,b�M�)Jp.!`/t�\���&�6mQc���ʫF��$K��]� ��ƭV|]{V�ffmc��l-1�e�`��TT"L����A��Q'��E�N1����ybǛ<L�����ҳW����0�xN��7����O�(�#9��;�)xW���1�uQ<�c7R�b2�&�86y�o=6\Rd�/��K@��sg#I��b0���ϐ���� ��/f����C��<y�\Sk��8��
�������0Dˬ�lr��`�u�#�g��A�}ޚ��h� ٢�I%Ѩ'R�t�g�ɍ�e���lWY����mɷ9����q_�N�~'�	�ʋ���֋S��S�m\���ܳ�n���q6�,6ga��$ʠ���n��'��BV+���-c,��|Nt#k�ѷX��ѩ�?���������J��!H�8�Z�w���+�G`/�?o�W��̈́�_�I��dW�>��i��;ي�s�t��/�}◂��;Yh�ө���sr�/���3�;���La*?L�V�߁�u���GSUmu����)����^~�IGDcY��(|�5�F|
p�i���a�t���׫pt.c��{�)�	��5v
���J����+e|����|��',bl�`��dc�q�Z-�����ķV|k� xfy�*�lD��|093>���%n��oƓG��� 1�b��#L!&0�DK��E���dF Y�9&��8WC�F�����҄���Dփѹ3���Ҏ ��t /�����'�	x� fZ�9P��P�4�OL&���]�8�h���Y�����"�tR&e��Fj�X������E�'�?�0���j5T�<�<�U�3M,A�|� 6T�+[
�Ɋ>/�5x$��q��u�n<z��~,�t���q6��"�pB�4���ބ��Y�`�Z�]�h��EO�Ô��R�4\�&.���7Z�Nݢ����gm
�L�]�v�U��(^Z�#���yj�g��:���i�[��g_�s#���3f��Q�D4\�"A���)��R�?0e��*ŋyW ���\�\P�O���0��-RV����c����}d�b"���6�c+�ƥc�po�������wjT�'v�XA��b���䇻tG�'s���qSf?ki��7��Wq�źb��\�Z�6���B���f�������p��(�h��,w�Z����U�8�&%a�%I�������K����ue�eML��{�R���V榏�
?E ����>TTEŽ�ر��$ "��ќU�¢P1����\xO[̡������J:�vE%z������aS��$�4h�=���o���{�˗�g��\�ܚH�G���$a�d���*�UƱbV��p�E}~TB�h��7�F����͝PR���4�>ՆR�:s��1CC[2���3y �K(��D@сw5�V�iP�ƫ���Zh�ؤ�1���k�+������l7�ه�,�$��$6�&����F �.N��R$Y����5�"���t'�}��l����ڠ���@`��XlxVHYEB    fa00    1340�w��Տ� ViA����Z��X��#84c�:b�m�`Qc�v��v`Wm�;��/i���=�z΂h�@��1�cDU�����;~l>��q��}�|=f�ѝ�U_��x����,Z����NQ�Q�|n1	#��J}+�j�]Dqu�g����1�J�����g��?;�21k�l�\�[�Qt�f���E�q�lRN��ӑO�dE��=t ��-9�cwx��� �E@�Q�%��ؕ����yD݌���&y�7gÄm�bR�ET?F1���s�L���7[Z��KhqyW|�m�԰�.&�Fd�s������qC�w�����nLa/�s� �K.%fH�����*2w�Jm��t��J�-�`�-s,�)vmH>�G~�@�
��Di�끻Fۅ>+��h��>tْ����3,)���ն���G��AN��R������q��C����O���Zwe��`�b�FrIHP�F���V�E�) ����9�_U�D�_!���"@�8���X��Wb�D���m��4���f�f ��l�r�dsi ��}����i͔�� �r��@�T.dЩ�(��P�TZ�%�I��p]wSE���;��땾2ZkYQ�Zi6SjP����[��T?�L�#ݝ�$��s`(���Pb�?~�>j5K���쒅��ϑ��.Y�j�:����^a��~�4΍��7Hb���{6q�^U�<��DWwD
k�a�]r?�T�x�C�O{CZ�!2Ϗ.iVs���X���5��ʔ��/��-b& ���]s������jW^���c�dp�;�8;L>[�?b���S¤ �@�;2\���7,��RD�}�<u_�8Sy�7M��&�ϹA�<:w�@�b�Xt霼��ݟ��]�����<^���2&���;�s�C�UD͚����
�>zٽ|{cCR���jE��5A��C��w�~�9P�������'@/Y���u�k%U���g�Y�Q%9@�u#�ɕ���39���Gd�Y��f�Ҩ�%߯�)�E�эy�ۋ�4�����\���=�7ٹ]�v�1K��j�1�Ip��x}� ���=A�m&�v�A��$͠�~�.=�HWl@R�̲����<rN�������h6Ʋp?��(x�>���7�����"/�> <4=�w�و��Ð" ī����⻂-��6c�a}���[b�k�K�А�{��^�"vݍ���b�B釰��F��tN�� ׂ��Ր}�PsнL7v��T���h�Dw)��b>�T��,�}�����{-�'�gp�x?�� �L���)~��17G��f�E�-L��D,���
�p��Օ#������ӝ����
�D�7���Omr�#P��U��压ѹU���9���&���`��������9��/P���՚Ό�=�	7}Z�զ�D��9�zd�&^��{�(f�pdiYp
e���B�O��k� �s�߁�!^ �7�9���N� �n�p\֞����Yb[i��qN���lg�l�_Un�a��VG��.wx9BV��f4e����2�C�7�3M��b�|+w�F�	���1p���`-��}:�Og���J���'��/eK��.�-mF������P~�5�|�	;Y���J�ʙ^��k'?N�U�����LW�K.�d����r����y���RO�q�Aj��xm]V�2Pt~�:�ω�>�Xef�����ZxK΋��X5R��zV���Z�{��é-,�X�B�K����t���L/�o�N����.9>U�X�}Ne�o���D���/*��E��"�"���k��h7"[��I&c��5�����*Q��m�JE�-f�i@���QӐ�E3��ʮ�^qg/�P�^�?k��R�V%X�ʛ���ϼ\�-C
�3bs��.�3 �JՁ��8c])�;�P�!Uw0\N�
������Yc�G{����,+=�6+�<�t�a��E�qG��u
�S;����!�`�s��M���
2�k��Ò�2 F0>��f�Q-�~fuJ�����tEFjԁ�Q�F��Rx�4?r}1>
E�do���s$n5�-BE���&8q�e�=/2��㦉^	��.�K;d�$o��T�c�`��4���$w73� ���Cծh�J����S`U2>��6l
�AԞd�f�f�x{�w�u+P*
A����z3�]�$�iL�Ϳy�g{��
+H^j��v�4��`�Ӝhr=ؒ.�}'�[e����zto��ۢY��~���"���)*ڸ]&L~U�ز��B��iI4��C�2't!5nl��\�>^�F)�S��DIn�4TV����	���cFM�T�g�W�s�R�&yzRU��Q)-k�2ioǴ��s�x�?�k��I����EiZ��RE��}��P��Ǿ�o��(y�ݺS�!��=�<�x�-0Z;�4�̽�4��ӛ���[áa{[;������_i6���N��a?d�F�n3�����&N��)�Pv�2dd4m�u��O���8�&ܵ"yr0���WB��5���Rp�د�ss	>���V��%�� A��\�Gϒ�!:�9@'/�ò)�vO���^�u ��["n���B�K�tX6�QF�0}_���t.3"���
�V9�L�R��$߀�O�`7�b������S#+d�l��{"��=� �X�PU������~bm����Z-ωq,�b*��v�K��V�G��,���Z�p�+W�xʡ�@B���+��t�}�����s9�{����"UVA����<�q4���B��;�0�n�:��#x��a|���Q1��ܟ���~�*��l�އX�c~x,�5!���:t.�����\>�9v�/r{�<o�DW���W_���1�wb���awF:s-y��CguR`5�n�[�_����PZ�#0�~�k+��*�o�67�SC��G�����N³�?�S֩X�x��3�"�)�c�����x��a8=e����A0ʍaC�����'>���#�v� ���<�l���<v��� R��z� �D�O�I��!K����C$#'�Q~w|_��UsNT�:�4k��47��D��!W̓�I��ԝ��x��"���Ƞ�q�]�o6O�>���蔓}�-�Rd�v���Ɯ����s��T�$����z�������fB_�<����'�!v�9N�2X���[��o��_����S(dv �z��>��M�!���;\�L��X~R.�	[7F���Mڷ����ˋ6��b�"����b���(�t�����M�qI	�o�����."���Z3�yJ&
Ŗ(7�AI>�sY�Ϫw����t��V�����WW`j�����]��ÿ�?e9Zލ��c��BF�7y��ǡ673"�.R�c�����cH.R���İ'�(�H�%"(
�6��;c�`A�E���_eƓ
����T�.��-�&��u9S��ӫ
��#�e(d�o��M�Z3�D�\�j<���t�ÃY$�~Hy�P�aO��\Ǟ���r¹6�̑��nJ�HT���n��	D���_[�,e�΃X2Y'��Ɨs�d�Yء�8E�>�>gaS��mLZ�D��~9�|i��7��,z��ho�IU�t�L�i�� vGT�/���+[J6���Ӝ���=γf=n4�u����gT���M��?1,3�A����wOM#��r#Ɏ-8P�T���L��6Q+lK
4R��@��\f�,�F(��N����I57K ���uJ���敨KMƺO�F������e����J@�#w7|^J�����r§�ad����"�;��x\�OSʇ
�����|�a٤�e��!���m5{zt	P9�ݦ���$ ��$��1���JǴSz�w3�62��k&��@�C�k�3��7V��^�(�^�I�m��B��A��3Q�w]z�s+V���3f�6�������Z��f�m��§�����5��h����`}���hY"7�7`*�v��=�+�[��{M��1����{t��P��T
��j��>"�S/��^��
a��:���k]O& ~�u\�j����t2�����OU%����:A�{�yXᭂ��6�F�K̿�O�8���c�#fy@�����"��+{03�7�6�~���|3�nm�F�;�0a�Z_�j���O/g�A����dx�#�<*���=C�ZfhE�.b(��(A�p��_��Y��y�^�4YN���~�B�0��s��e���kћ���x):� ��݈����c�֔A4_6Lut�f���.�6ߗ�@�`J���e�z���<��&Ϧ�4��S�a'�
�0��u���aB��EpsC���c�M�]�g�"*ƣVD�lp|L>22�6����p*V���pg	��8�"D� l����V�Ju��GS߽�}+r���#�pI+����X��TH����:ґg��S�Եl������mJY�YZ�p�-��_	!(�ظR;��:�#9���/,-�A93D�rl�3I%`r��Ys���T��ƒ�⇂xm�\Q�T��Y�ܟ����H�7��N=_�>{�(�+1�*��㦓�_�{��S�xX8�nǳU<�*�Ά*����D�j�1n��.��Ƃܠ)Z��$4�qu���<|w���E´5 ��(��D{`�����²��7�p�xB;��]��0���L�<Kg��߇-��g 
,*��F���o;�-̼&��l����Ԡ}Q��"|�z֑�j��i&��,�$�o�����4�7g��i�;;�A��#�2���3���FRW�z�mi�lN�(?q��E�"̕XlxVHYEB      e7      a0��s�~Vf�~� '�w�\��4٥^�@����D������i������fQW�'�,��o���W��&Y+C}=eS�鹁�>�(�"�se4/^����<u��J:F�EL�fe��*i�E���h&����#��ܛ�f�O���7��?Ej&���ihl�!��nr