XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=`a�T��1B��5��I�J�@׺Jߓy\-A{2A8���କFG�2&4���4�1~�O���
�H��,��Ċ`�$��������M}ُ���sV�ƷKv�1����L����$��P��귥�*��t*��j�{�_����\n��I�֑�����8(�"+B<%�G0cY#�گpk�aݽ��m�
���>��3�K���߾xY�O�J~�^������]E���N�Xˈ/�x�$���Еu�V���m6V���Hqh-�����ܯ���N���O�K�TH���"�|��y�������b�/,�J��Wk_?�=t,2x�@T
L��>w��C*�g͐~e�(�WnvR80�yh�⁖q���b��q`�l3���0٨��R���fp䇏���o�F��g;�TA8L�}��H�m㟗���ٍ8Ho�����?yZ��7,4͜���.fR�.�����PyP�E֬Z ��Y�a�,�lN�X����3���t0���E9�VWD"�N�؝�M�t�h����珶��C�4��ȳ���lp���H$����%��aQB����Tr`�+P���ɁV�����
��4w�b�IƯ<�H|�~y�Z8EvG��o�9B9�~��rl؀FĹo7o�|�XW�����*[��p�q�6y�Q`�\1�?�n��%����J�>��ڒ��ܣ�j�u�$�#�{�c�^�TV�Zg�T_F���r�^�Q.�{�1�t"o=�!XlxVHYEB    fa00    2020U ��y�{��kŽXy�&�a3VU�D���GRV'��ޞr�&��B-�`C�l�J%@6_?��n��$O88 �)N�\nM�Ɇ�����Y�K`�IkP�;F�:��m�gVeq����
P@�M[�z
��Rt�q�+�1(�'�".a6#4�Id�8����?�1�C��`�V��M�/x���ߨ�����&+�����hIEٚB�b��6f_5'����e��������lr(��Ee�[Xp���5�>p2)C�Fҧ@��%�2�%��go����E �U=��u�3	�]��=�'#��k��+)6ՒVYm.^���v��'{�~��^k�Z���f�m�Q1AJs{E�_u�J@}Z�s]7G��U�S��}�����ڎ�#��z�i��)��ڐA0sǗP�oK�	i<��=+x�C~���9]��B�1���Ipv�Vj����}�����2�Ş�B�ِ�lM�V��g{�����G�6�d�ū�b��C�e�'����{?_@*���ߠ�~Iі)I[�7���.�݋ϗ��]���u� ��&%��Z��D����EI������t3�Q�U��
�%�,���K�!�d�\Pv�?�w��3��Hx'���;�N�h{|��Y[���m킸�_�z�c�îg���}m���/�"���X+d��G������YvB���~e��U�Wƈ��"^���KnC�1c�1L�Qf�Ļ�^X�RK��U�Ye�E��'���m)�({�v�MZI��$�C�$���<ev�h;m��[��.V9�l��A2�BN�C)�k�l� �nϬÉ�6���E*����l	��{Z�1�਍H��%PT�?7�G��!��),"���z�c��6�����Ƌ���L����7,��<RJ�4r%ڥG�R[ι{Q��S��W�B;i՚��k4� 7�H@w�ܰ��x\��I����W�U��P_��*2T|��B�v��B֕UĒ��N�Ǫ+�'���~���?���.R�Y�]%q#�U����J�̰ng!��e��C�e���C�kT���-H��y��߈�!��B~��i�y*�8;�z��s���d�e�s5���F� U�0
�ؓ���)�۹IN�|/�\6*;�Ƹ�o�%ǚ�9�sl�����Q��ȭ➤F"�&�¹V��!�)����G{`|$�Q0�kN\�t-JX<0�.�õE��v�:B�IC�JI���k��A�ҭ���T�\]��M�X��n�0�{Ǒ�z
P��.�����WLb��<3�w.���EZ|$s�b���HdS!h�q���,��G�ob�n8v�P�!���K��{VҒѣH� �����O�h|ƪmt�,_)�X�(�k��c�%i��n��1��Ӻ���7}&v�Y����&l1Z��T{��@H�#JH�����z�(���f1�ؑP����t�n��[>3�5nB�א[��׫���
�^ko��h���~I�8F)뉒-kD_�>�����Ï��k���{êl���Eٗi��9�9��vƁ��<;_Zib��SU Lw�����M�eM ֫%���$TP��髡�]eVAG�P�� �AB�Qg�2�,���8����=�|���'���=�l'AW���*���Yey��d�L� y�/�4g���
�\8c������ ���[ ��"����BI�8���YQ����ި8�\t�,KO�>c����\�͇�#\���y�7$4b�2�CEl��A`��D�ĺ�
Z�2��S���q8����|�7�,�$JG���X&꼖Vf�H[ˎ�z���!s��U���V��e�c�0Ӭ�����]≀OlE�!`I
"����*�_�pq��7;C��Hۛ�9�ߒ�!z�lҖ �L������.�� ��Q[ʋ�Rٯ�Z� f����"���B~V�g��(����+6TA�s�G�M�N,l�����w���}*�Á�����jKPt�%�=AE$8�����|όrn:��nS@���^Z���_%��,?mJ��-19#��CRSU������u�[��į5�/.�^�j��s��F�#Xl!\v����i�4cŵH�������5ǵ~��45_y/���2a0^�V����|c)�����Lqɵq��r�?�=�qVV"��"����a�eUc	�<Vehl�-�� ���ke�>�G��~���a���=�J��b�Ea�*�5l��	@���&l���c���+A@*�}E�I�\���m�"�qDKU *�R����T��`.1�yS�7E%䦓a4*KA]ݻ��9�JzS�rѸ>:��?c�t�\���������_����-F�זH��uv@�w6�ZSw��+1g6���q
<*���F^t�0�h�����3�FQQQ=eùR/`
ant��Q�D����j0K��(r���y/p���J�;j�1����������<��nT��}g���6}�;�_: N��X����,�4�0w�R�t#4���x�!]�Z-�h�5�%n�:
h�%�i]��B�G�-{5$����'��7X�he=������m>������}���ҫP8���W��11�v��#cJ6G�MBC�/ȎD�O��P�:b��w�n��f��G���cm�vn	��(}EU�B8��zDq{����?��F�i'is�2,�^��~
aQ�c\ޛ�-x�!�6߽��	cv�\Ґ|��w4	�pU��@?/ɳM��%� m���������Ij��NJ5;[+��������������t��te����s&ٯX�N�6jbS��g�����x���cP�Q���d��t�,8��>�A�{��/��d8PF(=!�V�-���^m�ðS��XrV��֨�
RD",>�_%�����9L��p��v8+D��7b9�I}�~6�X���Z�Z��Y0� ����R��H w����ýJ�(�'p�Y�7�%;���� :��
zO��^�p̈́�Q@��;�~#y9�O�1X��$1Y0�p���O�6(r�cp*d�Y>�>?9�%ZzE���u��T�*�A�p{g�����`� 
�P���C�v�b���1���=$�Eb.���P���$C����QUw̋�d��]�����{_z�D>V|ţ!n�o���ygED�:6�J,�s\�C�O�����Xj��e�*��U���
/�1�@�����}�{����B*֢�a-p��b�:�4)���zy��Kv�+��^Mq?C�a3
�Ϳ=�<on
� ��L���c1e�W�O�X���6}��ez3��K���\�\(���~+-���G=���&fE+t�Dz6� ���&������t�����ɩ��QrJ���i8u��Y��74��̎@�h��8���,���b��|���bn2�x^�i�����9!��+�9�!a�\_��x��5�����xלW��|�o�]���[ �BR���OV5,:y�J�tI���#
X �G�\�+;�f�+���\#�O	�:e-��Z'Mq@F!7��,��z�zXV�t#��,�d����-�+�8l�ݪ�@
�]`~��ϓn�c��+ђ��*|;�G�tk����i�XFC��̹�V���}m�)��1?�����d�u��ڟT~]#ͱzI�֚5̾v�h�i���N}�w�(�����${�ew�+�4�ҡ��χK���Ļ����g��0�����b�fW�0�xI��L�ۗb���G�86H��f�����vodn�����i�׍Y��nH�C/�p?�����'�m�L1�_h���;�<s�J����iQ+����Z����ġ�y���ѣ�A8;�8���Y�1���t�u&�'�zO,�| �-�=V
 ���3�x��"�wo���/��&�����=B�g��(���i���}Qx{,��:ږg*�/� ���p����3�l.Y?{?MWA��7������R�pItGE�(�Ǒ?������)A�\�)z���s�ܮ�@��ݕ�<Q�]_h}F�sBν�����G)��t�Z4�����)-���� n2KC�@a�ME=sfw����Cе&�8Z��y/ۄ����xh�
W�^{O<��>%���]�̞�M��#	�$�ʂ�����L,ǈ�������^T.��y�Rwb��h|�!�e��M��]��/'��o�Wq
�#����.��=� eea��R%~{�4�ZK0<�A���� $fo���@=������'L�����HZ�r�]��4�+���|��Z� �_��Ɖ�|/S��j^x��sC�VAc�V�Ca����U��
��u�0Ij��8W��@Y�U)��)	Z ��(�Aw'���Q�}�4�%�j <�����-��\y�ߤ�Q���(����<�pEvl�����{2U�.�w�	nN��N��-�^ު;*�9����w5'n��})��#��̿"�$[O�%�l*�N���m=�����γ������Vf�c�7�m���r���k�gUOŃ�/�|��]��IZW�~ڢ(c��-�H���A0�4��w��:�﨔��s�Uh����k�N��}���:W?��8�Ħ����Pa�ZH�Q@��^l-b�]"q0�}�������6^Z��a�N7g��ʢ��<�)r�=�����&��N0(�f��ࠜB�� ���I-���o{�Ul�9���n�S�Guz��ZT�I�.��7$s̑��#W/��|S\�d����&�խx�_8�-�I�n+
w��2�Va�����zV���kO��k���qE�l苨~�Zz��݄CALɤ�����©���%&�JIXߪ�Y
m��9��-C�+�{>5$�4������Z�P�� (�$O�IG�v��W�a
Nu�L����e�\�`DS���4U�M�9��R����%����DFY�~�{�f* ب�c�#�rvn��7jc�/�oa�5����Inj+.��I�3����l��F�Bei@&"^�L�u!MG�Ey�_�U�֖���M�Q
q� �w4���S�R�]����V��P�@����i~�5���w?�Pт��m$5���`qe��#R�cc)y(��<Qa�?B)�.Ӛ���]�k 3en��Cn�����F�1ȫ՗�<�^��y�w$D���ǲc�:���w)SGlr��B�%va�7ٶû�k
���� �\㧌]�#(��W6;�t�qRl�۽@0D��4#!$�&c@��` �q#9�c��ҝ3��/��T=K������:�htn#�3k3[�h�s�{(u��Sy�,�	�5� Ͷ�b�~�	C#M�,X��)��j0¤W��i�>��#+����(�W�I�Ts�1I
E=٭~R⹮�h�c�%9ilA�]�SZA_Ud��=w���sv/����0^Ӳ���#�/�Uǭ��#:��7Z�1��:!��+l��Cl �|��z��!I�����\&o�l��=��l{UO'�5��<y�	Q	��7��z3q��h�Jf���Tp9��::��p��K�'8ٶ�da�ݦ7�=�QŴ�>�����Z>��JR�
�~�R�yp �Ո#Dh�z{Z��v���H��+�I�p�6�ߋr�~�@޹F�[�}�(���D�6�0#A�X�k` ���!�|vb����=��M��:xf�D��4;bǗ��0��L�O#�����#-~�j�*�ps�e蘟ϕo�(H$h��=�s̓�RB
Y��U<��v��;�Fkw̸`,�a�>�_����ę��-���ShN'd
�I�(�Y�4�C�[WMPMqS.}�>Sh;'��&��{]-^0�����9X�2�h�a�%^�e�L�O�F:��=��.:8�0G]c@[T������a��#���:��&�ZB����cάf�=+�m�vÉ���üM���SEnt��hXzpu���D���m\��:'R��)=�3��T��]�G�a?����y�~[� �����^��-v��st7���^X�Fwut�<0����������/�r($����-""�6}AJ)X�m�=�K�2� ��N�|6�J�����\ۀ����`���X��v"-��MQ8�?9���<fs���Zb��g��L�
t;P4�}~'�g��դ�i	�� �+����B,~ws���H�c�2R@v�c�)o�QI�c��H^�������q���B�@,g�i* ������\&�әٯ�+���1�ln ��"=~�%�r��<n�O|��+c�#��2�=d���R�:F�<��cʮ�S�j��+��Uj���>��7����#rg�[��D�7����#�~�g~�Y8���(��?[��Սu��X�y���kR��xc^��K�E�.�������K�>cOi�B����'O�W�N/)8O����,�ͳ4��Bk/�4�=��)�P:$��{�$t����^�u�I���W|���J��*�Oj~���!f���̒���e��D��U�H�{S*�X�	�~wtP��0L+�5w�.I~����ah�sр���p��n��-r0�WJs�ު��w��Mh��<�CGG�� �C����d��{�>����P�N�4�� _�������5t�E�J/���4�m䟩m��C���Kw�wt����R�0��7�S�0" �s�I��躰�{���[���w�EX6�V�7��r�0ս���u[��&c�4g�����"��o���t6�m*8��ZM�aa�'�M\]����L����\}��0v\��S34c3�C�(i*j���8��XR�ѳ��H5ߡ��5 �_�:+�&Zm?��d�*���J�(Sn�@ʹGu+�����w{U}
�J��@U�|}�&�>�}�릘���L�\&'깜@7a��}[�&�hK�/J�I�"q-�)Co���Y�\���C�؏p˿i�"���ˌ@bg���f�3�E-+R��?mm/m������_K�oN8(�>�s�K@����D��/�Qj�;`�P2�&b,�Zj�mtO�<A�i�
y#֥5���:H^}׬Uл�������3�?U�SI���a+FD���jmu8��A^�ĉЗ2jW5��}��g����	mٰ�
�{�G!�ntM;�&��%�O��l�>�;\�_��{� ��ie�%3�I$���}�~�t/�Fx��hS�|,�b�k�~�(��>=�J�G��� �gS
��l�u���8��Po�F�K��J��5?��O�.f{>b ���AZL��Q��t��9��$;8~%a��L��lL�f�*�'��"/�"A����Y���A�Oa��5R&7\�.��u\��.��_��� g-η�J#y˯S"5&��ُ��'%�)�a���Y ��T��:�|������{e/4�&­3�IX�e����q
F�=\Osu���T�l�w{K�b?�3^"8m��)�}��Mq�6ѭ�E�.�ܲ�gv]���F&��"zZً$>+\���W��O�VHj	~��� �A�P!Z_�iMqX݅�c �z?sVG���NF� #����5��Y�.�)`����/�	��\pnǝ�l�4&� ��:���`�)Ew��nM*D�RNd8A6USq����S��W�)�OI�0�����-��)Ts�z}�C�јd�r��.�U ������w`�J=v��/Z�/1����N�@q7�ihJ�Ds���o S��{�.4��Me��r�oz?y�)5-%�ZY����I8%r��rmzX���>.��n���0��C�W���mf�c��Vy�6��ѿ��L�޶g���'�r�Z�|�C�O����,}+�Z#�����}i��u݇9��
���{�j8�����Cʬ\/}��Q�st�K�ޕ2�M��5���|�0Ͼ���V��+���=P�q��k�dPX����!:�n���۳]	\���O�i���A�5�G��,��E@�&YzQ����yg���{��T(������u���;�]՚"�h7?}9�����Ϧ���%kͰ=�&��q��2,�܄`vgg�XlxVHYEB    cb82    12b0b<!/�3o�8��LX�|Z�fV���7�!>)Y�� �Y�e�U��7}N^
�-��~q�7c���e&�[`7#R|fDVM��L�G�5��e��g���Gq?�>�`(<u��ژ\�%zj�m��x���>`�.�9�:p��:2���d��Sԭ4J9V�g`�֛��c�v�������1�'4GȚ���j>�@�+�����T3ٓ��v�W�`9����}t�L��.g�,m�U+j��a}oĂ��q[S����/��A0.����ܛd<��K��X<I篼����ۊ㹝�௬�����0��ح�q�:B�'[v%g�#\����\ua��ؔ_0�����q��68�Vp�_�F$a
����%qל���"�EHl�9�"X�m�B[�!���9z�hh�v3�K�(m�:
 ��m
��_SR� �� ���V�8m�N��+��r�{��z�K8�S�	~)�%��#���Х6%�����+���^J��q%��;n[̅�.�0�.��c�{��l��O�W2�Q��H,�B�ٺC^�E	"5�ntd��~S0�bz4~ON0/Hx��]�E���ѹ��������p�m�5�־^c�K��F��FQ�_D8���vQ���E	p�ຈV�$�\u�x����Y7���CL�V[��4�Q�/�LX0�U�q]�<闓o��3�Ds�a[I���F\
��N��ʩBʦbE�(S�)󡪺f�.��ݕWG������=��ޤ��������-}��* �2��PIP�b�g.�E��dT��FH��TϮ��}Qk��M���A�������p� ��6cu��^�7�����y�.�}�-�c]��/��xͲ@��;�tNL���!O���S%�h�8-^wh:pr.��AO3|i'�����d)k��{w���V��D��7g�E�~�o$%��D� �?� 	�>�W�3)��~KBR9f(��EܖP��Xs�˩�WMn��7w�:�?8R���CFbj%��JO'R�6��>��$�y\Ӳ�"���0����
s�ԏO=Zh�#ί'z� ��خ�0Q⽝_M�<?n���˘ZGϰ��fy�U�a�Ԩc�b�y��8��H��G���yt�u����2�!;�����`� ���*��A�Ǟ�B��$iq�ۇ������?�@2�>�z�e�t܌3׻��N	�ζz���M�v��UZ���xr�}����T���%}���+Z�P8{Ƞ�K�M����W7fĹ<�Hob���!�^{����d��Z�2SG�W�	xW)/dޕ+!W�����bT��U�WaĶ���Щ�"z ؘDK![�ѡ�z��.�u��'X�M;O�I%U�6��L��fG ö�s�q�T���Kꌦ=.�in�7��Ḟq��7B�������ťBd�8E��X�TXB��N��w��s����m+2��ƮjQ��Sh��m��b��^(��(H��U񅄗���P�U�u8�ۘ����:�����*��%"��_�t	�Q[����c���+�*�uC�D9U����+U�Ї� �Hd������\rUq��/u�y����G8Z�x$������v��m�ken��NX�VzMΗT�[V2�c=����3z���J?w}PI� )I+Z_��k����@�7�!�,{t%�+%Y�8�����@m.�pZK���VS=��z�����~�'���|�'�-\�7P���P�(y�ֽ1>�L�
�JW3d�|�P��6���l�y��8t� \Q�/�$�K�����t�W��w[j �7�Ù�Wy�ϖ\��b�sj�*~&��ɲ�$?�S$#�%����hg:����
�8N�^��^\�����7�ڴL ����^��>v[�/L�ٙŬ/��}��z&N8��PRa�3ғ`~@�Z��qh�Ӂ������ '�|��H4�ԛ �c��s�3bQ�YE�����/��[�M>��°'��˹BaV��w�Gn>�Â�E �sEj#
Wj��̺�I�2:�D���3Uv&7�$�L�K����,���$�u���/�}�PLu"�����?'Uw ��=�nV�O�W�Ou�M�u1_�>[���$_9냽LHH�҄t�L�����FR���WnVr�v�Sk潅6}��J�Z��n�K��e'2�Z�Z^p�N��@8��{�"-�-�Y${�D���� ���+�tv��MW��ɯ��Fn]�@�o�������xy�
3}CS[`C����R���T��dmɭ2����O�A��O/>[��o"����䑛�QX@��N�W~���B/�����LPϸl�NL�iXV!�l��=,o�N�=e�&��R��
 ��W}��/
W�u�W�"I4q�mUcY�"Yn����smp2��XA�	��d�_j� �M�v�[Ni����K��`[�穒׭�`����퉆�����\OS��g@r�,��x�2��(��&���m.��*f]�� E
H+���1�<뾩��T��,Ư����iO%8�O�;m�����2�m�.�z�4uJ?�^x�B����j�58�s�Q�vM�OfK��MMUߩ8΄����&=�F�e��F�:I�7�z�Ǖ�&Uy�� ��<ݤ-2�{�]�֩��R����İ��1lg�R%�s�z�ȵ�xsn&q���t��[�;���S~��5R��0�-t=�`�[p|/��gW e�g�Vҋ[��dm>�I����B >�5>~����0�˲"䀢o�;��D^����|�a�ǂ�2o��c�C��I��}p��A_���C��ׇ����}��(a w(2�	�1k��`�˺�}�w�/��͉W�K�禛E5��./A9|8���K�D����i��J�{}3�&/���cm	}Og�ʕ���װ��7���2y��#���a��p�]���ry�a2��-Y�Uں3t�TZ�h��H��ޠ�y@�z��𝮘+J�Q��}���k��;g�~1�u�G���0�"�,t/{��i��H��e�|�,�/m�������Q�YCY��*ƶV�|+��Qj2dp�� ��.�>�,�נO��~pD�G Mk+>�	lh�n���+gB��U�� ��rƒ
�^yjTr3?�ݝ*�:�-}��'���ٕ��/Tj�ᾐ�34-�������ƲRP���
��:z��y'��=�'�^6�D<�K[���Fe>���:��9�(�!�*K<��˫k���/i��M#���A��N��Zкch
�Ըۘ"4�	{�_�k�{���a]��C���Q.���bh�`��Q���1}�ws����ؐfP���.K}�=al�P2F����$��G���+F-&��J�ѻ����$��"��w���W�ө�7�z$u	�e�s��2�)QT�Crwʆ7	�=�_ s�S���U�}�o����}2����Nȷ�v��@�:�#�7��F>�A��;��+,p(���D'� �Hђ@��<y����v�I�Ч��7`�B�j��_F��)��R�6��P̓���U�&"�K/�B�\��'�I_]�B ࠲��M�ڂG2�o-�s�H��D��XC�`_�����{?h�Jk]y��2�������8y�և*�Y�0M�~�a�ЈW��?u�ZA�R�y7�9�}.�&q¶
[����gŃ9�k}�]�&�\ɨ��;��HV�N'Ç�v�x�!�c�����t��Wީ���~Վ|�
]���颀�zt�C?p#%�Ð�3-3�$Wh�9���ҿ�ֶwy���啮�Y.D��ֽ�d��K�iL=������d+���:T���/�̎4̬��������?}�J�5�������*�ޖp��n��F� "��'h:�f��̙h]��O���\�n���|w�R1Adx��*�NY�ˣ�'�w�a�|���H���e�v4��իe�~x��g�'d��e�HDպ(�"UW���\vr,���o�
��s��\B����k�fP�K�������<�Ҍ��;����3佚�,飮g�'�:)���S�ba�]Ϥr�	a�	��1BU�Q1F_�2(»����.hN&{xɜP�D�g�b��r��bd�	�e�:�"�81���.n�E�I��%�w�+�;-�*���4�?6ICyߴ�����7��Ų�܎P�O��������0u!���r��Xz�٤qu�*��:�z�%#+�z��wTC�-����9�Ol$���$5{��YSL���挳�"E'-㒩�Tb����C�D�VV �Hj�~@����J�p���isx�	�����N��N c��S����v�:g��XuǙX`p�,��n3X$6 L#uU�`�N�$��B�}�`�h���������Ĳ��2�@�_���b���e�.9%�r^N����]��B��XΕz�d���� �B��/��Lj~
]�b��3���B(e�	�x�P1Ӱ� (��P"��vQ&8����Ɓ�d�h}�m2���k�� ��Pf|\�D�q��AR�ަ���e�4���M�1 CZI���e:#�<k�)0��,��������/�pʇ���&'��ȅfS5�D����,j4�x@�����s��.�A��b����M�:θ\X�#N��!4ߣ�7r�hW$<�P4�<��k1 �/'����<�;e��P�� �c
�,������$0:�	%�`���X�����[�k��Ø{�l�4�R|�$����WM?���]|�h