XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W^��
�^j��h$*��_��(��g��w$�� �H��ň:�3��(�'˫��I)�B_�K�^c��-7t����GR*<�ged;�<`M�&�@��?
��BH�c]�B�|�v#����Z�%�(�M��[�� �foW<�P݅R�������D��e�3���Ѭ��+"a �άp��|�F:T�LO�Ɩ��A�C�g� E�����D�j�o,�Y\F�.��E{\�ֶ�Xz�r[L���΢ ���f9�fw�)�H �w3��EA�t��8���`s��[�Զ�#<�@�wom=@dq���E�A���s�9�]w��_���n`���2���;|�����Q��������,hp�R��/�z�h$"8>h�u;�D�6$������:�~�2�J=����i�V��GtM>2��!�&�M�� �L�ہ�̦�ϘǱ$���9�@��V�WC���g�\��Yt��O@��)[
4���x;��_���YP������`�:ĥ_A�x���Ӗ� ܬ���T�P��c(ٕ��A	�ioQ;6��9��[�l�]�l���p���^�w�MAA�id�4���Gs���Wm��,�o�(+�ǾA�z>u^p�<8��h���hC���Py�9,sO�&�cs92�a��Ѻ��Fф^��4ݻ.�{��F]��/,ݚdH��!���ԇ�Z��#7g����"�p�@1��K$��&_��r�/4�0��������菆�x�0+kXlxVHYEB    162c     850k~�/ch���uk�LP���$%r�(,�W��9���n���*hc�\�Is�*����8�.	�@q�J���P��ϛ݀�1WH�(FO��2������Y�8�� �j~�S�T�Nո���ކ�s۰�3����� �1���n��k�"��c��yt��0;�tx�Z#B�o�B�s��@^3�)X�؈ݩ�)�"2b���uG�K�W����S�Ԛt��t�&��L�{Tzq7�?�t�z{U!u��C�� �/�	ŏ,{�cm��ʋ��Z��@�Y-�B 3芎ZET:��o�\�v�X�V��Fx�^ ����)� ��`�U�(x.�������p��O8���T���dƢ806�v�Je��3t<�P��2Rq��a��~,������X���@벮#c�{������Oz��Jώ�ih�$��k�	�JM���w�(�2�zh�3<�)�E1�t�����2�(t��"�� ���m\v����K�(������R��ÿC���
{ �f��B������7� \w�b��=��s�����5��~�l9*6As�.���3��l�y��1??y�*ߛ���Z��?��5�迳���l���u�KݹqH�4�@0 ��B��QhX�����!#�����α�a��\��`F�z�*��9h����jW݁ ���n�u���@(v���kx)�&�K���EwF��B�ʥ���oq��)��ʼ���xzJv�>!?����}LF�z�$�@�\H�d�&��2gu�b��e�ag0�d���k�"��+�;�����@���6F������6X$�
2X���e�5x�s7H�8�t2�`.fXPr1��y �ѺY�{˵����l#��'<�+g�(�.ML}T�D��@�PO��&��&{�y�Dʒ����̚�4�!��q��� 	���,Ε�;'|��Y�"�����n���Gӊ�4gh�!�ZU�a�k=���2��tY���k薻��1����y�`�ƧN�
��0`#
�ٿ`4�n�ś�Կ��%rNN^��9}��?`��{�N�=o���\a�$Y��(D=,�k���i�ۇ�}�	\�|K/�G�kD&5����mz���+������K�'�j�K�Q�U�,�MnZ�/6���2 H�t<?po����g+�R
nI!��X콜���6��S))��J�T0E�ﶚG�Ц�tc�^0��Hշ )��O�L`���[+�u���2��v�S*0�o���z.#��Vnݯj��6+���Ÿ_�@�j�	E\�a%��ԫ,���~�]�J�r�$��K�ߏ�93��Tz�m�,D8��g�8�?]Lѱ�AVC,j��p�R�.3�c+��\����;����fLQQ�?���Q>*a5��rd�;�P��u���"G`{�����aBK�$�	�p�;�����Q�����֍���c��l���0�	r�E�������LSH�����g~��kW<7�\���e�M��A���0[O奿��x;$r��g��ܡ)UԳ�/��0�L�vf�@�6� �Q�"�^B��恻D�a��&\P�([�}`I�Fkb����8�3V���
�ց|뒕U��q�rv�=�l@^���)���Je��g{�����x+�����&�F�t�n�S��<��[cX9K��Ɯ%:�7��p��fͱQb(J��ax�9�V��F��m��6�^�p'�U��:�'���.��ȎD]fJ��Ukn��A���I�� �~��u~I.;oH�:�u�\�aR���oZޛB��UT!�j��$`*�1�^�O64c� pw�=������?&�+3����>��ʡ�K�kƐ́�	�E�4���"er`�f&h�ү0���/^�rȘ�z�KO@�z!Gb,՞m�ҿI��k�:��N��mX�}ZD�F��fN�?Wۚֹ\�wNH�4��-�}�bE����2��\0L��>��}�i� �� c�~�؜�QG��n���H?����9��i�K�p��O�PA�.OwB��L�]�3k�iՕsY�6��U�ޒt��j�-ˢ�����~���Z*��=%IQ�s�W/n;s