XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��sWT�6�N����^\I��=jk��ܘ~@N��Z~��Ӣ�G"?�F���(e��Q9��]T䒬���_ ���޲�9�	G�nk�IQ�@�/9��6B�e��o� %��Ky��mJ�c�|+s���l���%g������B/ł4[y���6Jub��,Ǐ����Z�
��F3*=v3�����0�Il�|�X��ݛq��Ɖ �mIܰ��O�s��������qF"��L��)ݲ~���w�N��*۞�h|V�Qk%�GD�F�_�r�#�A?�`O�S暳'Ԯ�Qf����wLz{��BAʳ��율��k��j��(E��Xۖ�3!�?���V��f���
F����J�T��>5���׃�����h���	\sۀ��2��j��	k��XP|c�͋�n��U�5R�I$">V��ð��q���4��HF�\��od&cs)�	�%^��1����$��[Nn�𨻢"=G�6���)��mð��_�����v�$���
O�4l� �}W��N��6�����kCh�t;�R5�mˣ)��k�1gAF5��R�t��X2�F]e����2�A���T)��E�D�Z�˱��.6�g#.��$~9{�HU�+Z�MME��ib�

Ɣ@��2�?/Q=T%y	惇�-�:%�JXl #�O����M���ї�̕�A�A��{�6w��O^��d�{�4>������G�.����+j+[����XlxVHYEB    4089     e40��S��i�9�MoX~�����x���sz'�#�3J ٬Q`�/��A�t���-��*�I��_	PR���y�RS��_
�2"��,L��=£�D�������mG#��Rw93�|���"*u�a�6Q@�Q���m'xл9�Gk�)���n�A�0.����	�=�j
���6��U�v�:qЃ�vɄ��;õ���F@��Z��e�?�^3�1�@��J����:�����B�@F�����'dKzc�-��F�td�'��nz9_T��S��j%K`�2$����.s��P{�z $򎠝Ў����NO&
����+S�"���֕�����&I#|�xN�v
��v9�e0��_���Z�l�j��2���`�j�$�u$�6�� ��y�vb�W�\���a&Ip����36�N��BsΧ�o&�(�;o�K
2�ĝ�_U�^�?1�Z��C��%�+ͱ-��%�U��҇ɀ�AP���q����Y�n�
a�Q[���wq�xSy���H��:�efl�<���-b��޷�y\T�&pIwn� }�2�O'��}�����\��u@��.q��Mc-��԰�w�?������	qj��(k	R�_�r$dp�D�{91?
2��J��nx/�!�A�Ȼ�1e_g��_��T�F����%�(�	q~�hw��`�s�X�֎��j¶��D݄����vnwT���G��Eq|ap���a~%).A)!�
wc&k���{:�O%R��w���>�?�q4�p0�;5ւ�H\�7EC��4��+T�X��.�V&(d�~2mXK���KS�$���ӂ��B)���cQ)���ǜUˈ�@�w367��wsPBv\@{���6�� G���p�.;q���ܮ<(D��K��x�?��h	�� [�wz�z�:(/�pÖ�nY/
j����&��H�KS1az�0mX*HE�@¢���m�}�̏ �XB�C���$
�薂��=	���A=e)_0>�q����C�z�sh�d���X5�ھ(u9M��:���s<I#�ݓ�}^o���L6)x#҇èHs�}hP�i����:�RM�հ˓�'�
���ɂ3���%�8���Z���؈��̮�r��XˡJ�B��Z�y��E �K-޳H�"3�<6v�|Ve���a�' �w�J*Ϩ$[�aR��"�S��.;�Ŀ���(���/!}�l�I�o'V;2�Y=�I��d�{����|�d¹�E�$M�|���gt=�`��z��9Н	J�훓�0:
=�<�uHπh+�:�\s�� �ai"q��`��8E	�fB�L�:�>�ڌ���:��V����2hJ/%kh,�y~\�Y"L�f�����`sl;`WԮw���~�.�K�2R1��<F��4'����s�t�b&�l3�6��k +�}�&|n��J����� �ad�~���>	(<���I��,r��̛q�%E�e{s�;g���I�m��R�Q�o2����U��9�1��f��C�ڟ6E8�@/��[a~O4>E����Ơ�X�M4)��R��FBv~V�;lu��1�jwO�DJ�EL%P�1��6�d6GR`���,�Q%�����(,�/�Ѻ+5'�u�}xz�� �Pov��_�,�����|�5����#�dO��4�x<:G�`������&Ӣ��b���̀A~�É���{r����O�u��[���d��%��በTs�Ȍ�ŷ�x�����=(-,>+<���4���
r�YȐ����RyQ�����i��|B������^�����T�[/K���V�vqӛ�ϴT7�]�jRn���DF�ʼ�Ƿ^����Ɠ8+SKL���hW0�N@W���ʗ>E!��xU.���yV�~Cm��V���������c��s�M2���æ�e�%�?k�J��8;�����K��|���L��~�A���^�/��][IO�2����aQ��v>2I����]���eH~$��x<M���&<�A��.R?�7L�Lr�+�|G�l�H�l�a�Ŧ��6�k�p �k%���|!w;;�u���Z�$"�	�ρ�v
��$FI�W�P.�0%��$é���\���M�M����O�^M��������B,n��m7�R���t� A2PNa�ORؒ/h��V���w�~�E	����X�[�]V�����8�X�[�y{��+85��`�L ���� ���:<���)y�rz���u��@f���J���fd�v^zW�~L��Pn�vu��ـ��PQ�\����o?�¹|�boQ��j5�k����u�f�9-
��&_��r��u�u�9�!���
8.��|�^Rj��E�[��?	r:{��èzCƌц����h �Z�n�YĠ%A���~��]R�'B�0؁_��z�5ei8���a�����Eɻnvj����w�Y{��E���		�Z��Q<����@�:|$�u ۈRQl�W��<'���1�����_�wi��&�-כ
���Rk�n F/*�'pE�8s�VXҖ�k�Ke�����%K���MzM)�S�Eo`��w���Ym�:s[�n�D�(>P�������A���F��wV�"X��r��j���P����0�Z6\�H'�]5�X��Cr���i�í���F ~��-*���ʸ��=�` ��(YS�dM�J+;�/,�ᚖ�tV,�ACr?n� �����7PU��� �iװp���!�
�P�~K�`�̚����Y�Xj7M��+t9
ע��%�K?�U8N�8;�J�����^�S!�N����3��$fy�� T���LȦl���w��nǢ�ӣS���
Ց[x	U��U�45��)1� \��k��?2�����y)5�_�����,��Ok@�Z�-n����E��|�{sFh�
�p����2HFL>�*���^W��7���9\Nj!%3�ΰAz)m�c!�jq*K`���z u1`KT�K��'��w�YU"Ϩ��е#4�!�Q��ä+�f�'~���@����T���ԭw�����9믐�C��9��ϡ����ҍ��u��"���t�4`1���TL{���G�
�)��%� ֈ{2��;>I�PH�y>�;j&4}1�I�gPo�w��qL�$](���g�@��-��-�(�����4M�oe9���~#\$��,&a*��Z5ˈށb�c
_J�u��q)cI9�RF�Yv�c�|	��q�GY��ܶ�"�+n�3�<"l-F��b�*�"?���%�� ���Gz*��č�R��.\Ѯ���'`BX־�x-'��J�^�efg*�Uڹ�چ��o'�������z/B��Ѱ!�}�g��j��e����S �A�|��%p����b�ʭ�@����<�J�JF���G��&��F�Ӣ�z��E<��MLI�R��NB��
ejg7�?ʼ(����c��C���4�X�H�5oБz�n�2����>xt=Vq�uM�_.��ۅL��b�^�0P�^@���M�pt���L�"JJÏ�o>�r��/�!��L,�϶LŔ������n9�ǖ����EC7;�fyj��0���Y{c��k|����y��V�`R�&����K�_�V�}���t.a��cQ�