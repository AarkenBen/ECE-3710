XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Yh`r�ǵP�2�����7Ъ� D07@rW�*�n֍�?���uƻ�^�ڬES�yBןV�ɠ�E/ƐY���H}��D2�N;�i�i�c/&�u�͗\���]�qit��#��4�ԉ���N�g���OU����A��c��\���������\�Nn%.������h���to�����$�6 ���f�,7S�H'SS�P�v;�a���[�M�?9;BT�@��[�!�{�`½���wI�
wR_&�'7�6w������f���X��=.�ݾ���)֭�%�P$���(&JRf�z�ֽR�J�푈����"	�7��WBj<�����x����gK6��^������
0�D���4SYA�W���rvy�͸V7?�&J|��f�?����uK4�h���[!D��[�b�.>�ѵ���F�C>,p[���%������wD�ɝGI�;���+�*�%���$vYUl�f��\_G���x|e��70s��Y�%�b�?�h� 'o�����EP�����Q�R>S�1����5���9�(��a��b����/%{ԇ�!�}���v2ԳY;<%:�,&��n���l;��'q�"�����e�1ӑ����W���,
�=�����Vg��H�*���uGtRwt���5��Y(������I)��ז���&����Pp0�ݛ��K*�iA2��OڋfVJ���_=�oX�*�j_\�] [ϡT�
ހ��֧_ݥ�M���XlxVHYEB    fa00    2560�=(��-i�yR��=�YK2^�b�O���hlQ���D�Ul5ԏ)���qK]y�r�2BԓF�:(�w���� �W���uu��"���@�6���&�&\��^�t������C�}z&-�.�U!W1���^�|��'�CUI�s4N���I���x�?�~̰|LZ[�Q��3�����AG�S�$l�������Ϸ2dA��T�sq��ǳ]���)���x�P~�y�԰$6�&S���obmɍ(�9샑lv�z��3Qjd%�����rzԠ��f;Κ�N��@+ĸ�t�-'�͚������N;C��K][i�5��d��e�!↘J��Q�Հ-�஠W��Y�R�o˜���1Ql]�+�O�P6+i���ޏ		��a�h_i#���$	�����3^�Q%�N!%(?be��U�s��!S�+��`��2P޸R�5��+�]3�	f���[�+��	wE��~�u�D�Vs������v���f�Z�<Խ��WOw�+/�9��LS���u�$ Y��'[\=+�����`_��y���w憍:��V�w5C�������A�O���t\+�"kFm�~=�G�V�ߡ��s�Ȱ]cB�����dR���N#t.Բ^"w�&���ʜ�[�ao�cq� s�"�{K�cg��=9�֖ݰ˙��q�W�6�>��E˺Za�F�27}|�x��-R�z"z{��!}�DJ��U���F��ˈa����D'��#H-���t禑�;$�vپ3��_%�o��$6�HY�I�:|��M���}�\?���"Ry�nU������	%O��;"�6~<?��M Y���h�!k`FRCǕ ��XFd���s%�)37(���_�>}q����*�\������/|�|UO�D��;�FI����mwܻ�`��3��t�y��>,�Z�e��A�H�!D�Jc���:Q�D�B�L/���o��i���3��g�]���<F$u���������.��.����.�B��n�e�C�ܝ��c��p����p��x�Q$rG� �yВ���:g��ͩIP��<((�5�M�(T<u�*����|��0���;��wK.���qw;~E��k@?pZ����-�!z}���=/��[�?�$��ԕ�.�C�ʒ�`��r��S}zj�jC�}�W�b5�o`Sx+}�L���;�x���Ey��0�/�pv �?�ђ�e��'dr�s򑸬<r��ڈR�� �_/�
�C�W�$���9��/��M~ ���4���;K���|ÚxQX��3�_B������INn�r苝݁�Uc��+�h�`�z8cA�YOJX�|I��Mv@mM��Abxi�q%�����Ii�J;6�̓4�p�CF��gw�į��e��r��)�e�Ҙ�-�L�A�:�hMt�^�y���=�B}33�e>�F�S�"4��)�N����%_o�wA!1z�U�L<�1e%�߅5<�aX�)��=+#@����.ۥ!������R!"�s�(=pQ쁂K����>Ћ/%���P���D����1��@��E&�	��즗���9"w]E�ϒ�l��.��V�]M��DM)E(�	O��˞2�i�Y���=�����QT�b�(䅒� �u= Z�^ �3����z�S��w7���Og:��[G���~>.	��I��!� ))o�!�����%�|N��-���u����f2�0FŅ6���i��q��� �A*����X.�3q���k�U�������7]|�@5o�5�?��&B1%i�/ &�D���WC=e�%ѢDmw4��ەc�i���Ŵ �?8�N�9EƷ}MF��s����k�8<3&7�V�D�zˈ9Pߌ��.N�2j��?�����������j����5�6m2#�b�޲T�[Y<bo�z&zp�9��rU}�Ě=���}#-N�0q��W�In�h���4��
�4�F���<(p��-:s�W5����� �^���hSKL4�d�P
Т���T����BB1%ӷڇB8[�V�6l�5�+�Zw�(��@�� 1�Vh��U_���aut�a�U��"��~_7[%q�-��R4���-��f��Y\Q��]ܶU�����!�ٸY_�:d��W/����h�v��?o��בgK<yQ;Y�C&b%WG�a�P�!�v�})/�&�r�y�����H�s�y�DD -�f�䀝�NjHŐ��͒��}�+.�]}�e��3�X�3��ߓX�k�㵐��h���ܐj���K�#lJ�y��cv���y��CŚ��mw�k�lwGMk:P҅�L{*��e ��e��/ls!��EZ��&�t�n�|���3Gn?M��q�}��h��b��C4�WmQ>�Wb���I��o�D\�Q	N���Poɳ�2q-Sa���ʉj��3�hmY>u�x*]/K�(�G�ȲN\K �g[<]``��nE��Ef�>�6T�Xz��R�Q)�4�2f��F[u�ϩH]T����q�}���������\�U#�q��To�&�k�B'�u��ݢЅn�;{�Kbz`�,�i�� )J}UŁ���{�����5��نJ������t�!��[��)YC�o��q�_v�Ȩ/���D�	�K�~ևpj�2�XRm.UC�C��|�D#j�`
N�Qf7
�+���r��8|7�v�O.�ٴ P5L�bU�p%�#�l@S�������-��~S����0�J����-���-�~.��k�˕��/nx:~�i0 �'�eh�^z꼯Pj.8ڌ���(�����c�R��lj�n��{4�e@D�1��  �����L�m �h�θ�ƾA�.sv4�k{�æQ�
6� � �N�اAN[�����ҫ<�o�<�kv�<����&F{Knk�&m����Z����3�,��������+�3�dGj]�%�p�9��QQgS�����ڿY�dU�n�w�����Bs�dn`o��W������L;�-����u�H�=�J�V;�ԛ��嚎�*xiA*�N�Hbͼ���g|�,�eElr]7�OA����ҳ�s'��`FX�Y+��m1)R��j�qG�t�6���,"�)w�Z�r�VUaW�4��T̝ �~�3t8�ΓngQ�5�O�� �~���#��ġ�zZ"���׌��緜7ܘ��2[_}�������6�L����UAi*f�������a%��9/�(_���>efU��ݢ���@�1��V�X�4n-���(�k��lI���=|ՙ�@�D����ӥ*j�`��I��j^�W�{vDX{Y$)�ߴH�F#Ң��,r ��B��Ҥ�h���>%
z�S�`�5�.^����Қ��aBBz#�x�mD�e��-M.�*[U��\��˿��JThr�@��F%fR�V��l��w�p79x��wW��V��YU�0�7�׫I�XR8^ҟ�_Q{n�l��}� n [|Lkvx%����Mi?��� �`��v]�&A�^Wc�{f��A�����B8c�k@��*ߨ	�hr�ɂ���>)�~xM�K19��[N�Z�Ҥ�>!��ȳBZi�F��E�o\m��A"��>l�U@�#h��)��˼���o�_%eM��t��7n��`�_�����r�_+�U-�$�-�j�J�I��K�V� �Z���+�gJ��D��K�]�/����k�>mO��9h(�K^��v���
�]N�m��na}qQ����8�Ü�����~t�lu��P[ܰ6(�n�X3e�$*�4!�x��ХOL=�Ժ�C<d"�V��ʈ�T� p��ZK�z3�"Y�ua�K��V���	>�m�s��L�ē�'_J��<���}�_�	z&'��,����z�'�=p���(c�����9�Q
��B:Lg&�VQ��1�nY��rk��X�R�1Y`�3�'��S&��'�xI���4��_��}o���I����|}��y�S<�o%cQ�m*F@�4R@��.Q�k����	�r�j�+l����m��>f���7O*0����6u	�l�|iOׄ���Sl�a*x����H$[�t�m񞂽w�Ʊ4b�E�z-�;�O,y1j����P�>$a_�����4�:�RDk3nG`靓��
,���/+�1�5
V���י�:u̟�#�FA����zb��U��� kB�;�)��m�!WYr��-�CJo��BaxJ�|�Q�-/?��:2ǳ͖� ��@����6�xA1�2zդFܫl�c���V�K�=ڒ\��ѓ��G
�X�X@`�t�k�s�xڕV��/�����*�ju�<����3dLP�{hi~|�w�7�'#<!�UO��Qh<�Ac��]ܼߓ�A3j	UƠ�G����1MVW���:mH҆�5��I0�P���i�p�ಽ���qe�U��{�wT��5�z�bk�8l���1 'g�iw� zR,���G)��9�,�@ ����,�;�屐��U�)6�s�����$+c7� Q/1j�%Ѿ@�^:���\��Vn$Ո�h���z�84.ƀ*Ľ�}�D�$�!�����+�|-�ꂺ���u�vK��>�~g�������2J>Q�����4���l��.1ؿ%+��S�T ���B��S�n=���H2K(�<.^��y~glX��p^"��-��E�����r4F��!6���L����l�gA�v�?�"�s�����S�I�[��	n��a-	�(��PT�qk�ˆ-'H$\�(*Ç ���F�����l���&����ǐ����<:$bV�OP������jMˇ�ڇ���nW�Q�l�M�߿��t�WL S�u�Bs]���Z�FV�$R.�_�Vy�6~��<�W�9X���o�U�3����lOM'	'Y�T�R=����B�q�]��ui�:�Rч���w"�e[�,��*���t��&=��b�^��cРe�W]Y0���	We:ȑS�\o�\N'.�&E��Jl�pm�C�X�dd^#/q��<�s^;���笓�!�vb�#��1�,�P�{�S0������@���G�@���R�;�����H����W
3GUDU$�f]��� %B]p�x�T{��b �z���E��d���P8�QL$$�9������%#l|��NO�Q��t�=�#r5L!|̵rq$y��m^��¢K�[H}�1�38[zw%��#kW�l^� ;qNhAV��.�eUp�U�o�t��DCT�����8�kg��>@�&8��j�s?p��;��3�P�M�ͱ�tE��^E@�%����Eq3����%�<c�R٘���h!�_(4�ͼ���<�h4�y|ED�Tac�P�@�v�|=�[G=��L�O�$";��(4�d��h/XL�FѰ���{iE���~<���~�ލ��+`Ab#_7n���0�S��\���$9�t�輙���h�{�kٟ	�����w�zb��8l�]��~Kް�"֔��d�-��"pV���vƥ���?�!ܚr-R#\˺�a��iW�j\U[v	���}�V>�I((I9
�����FJm-	�� ]P�)���L]����׸QH�5��a%v�%����Ϝ��jʙ�a��ف�m��%= ��H�c��йT��������J�M�=���)��κ�
fy��Fo��\#f|~eZ��_C��]@m�Xu���5��t[� �'�i������,�&A�[{�l	9���������@cwAD^���s���p��k�'2�];⯨j���"� 7Դ_���D/!��1X�H�)`�F\Y#�I��}�i����5��H�(�t'bnl���YU��_�/�'&�|����q�8/R?���{.a �;�~h�=��|�W������3��5��S}���'�p=������1O�IZ� g#'̚k����J2Y�b�vJ|y�caiXE�`�k�pya<����o9*�����C��,
B����`W�Y��d�rTɓ�Βv��#l�%��7��/94M[j�D��3
:z+��T��f��.�':��������x����\ȕ�@�4ߨ2��M�9��Q��y$�p/[���Ύ`į ���|T��U˚�����H��(H6�	-����w�h��o�ݻҝ�/���X�9n>�V��Tܛ���K@6,��n�塑������%C�V�^�-E�.���No��G��-~��b�}dX�<����a����'"t�w�?���2�Q�O�����@~�o�c?�����n#%�y�
�K�z˘���c�q�`.�K��55��J�#���Z���R��&��U���E������>!^ie�u%L��_������"�w��w����>SL�j�w�)�H �,Fc�If^_= |�� B�#2|�>J��ɟ�I���K~�pH�b�w)��m���;|��O��^�l���dy�PI���i� ��%�r̨0>M�޳�(�R����Lqs��ř8TQ�2��Հ��N`%�8Ou��<#%t��&�'%��Z#��/>F�}�T����y�X��a����僲@��<�ط���'����]��-��ކ�F�__�$늑�Ӷ�U6{e�O��{B���O�]+sr�]� d�9r~ŬT����?�L�>7�v	Ȗ��C�~��:���-�'���+*�T�Ā7r��W�jC� 1[��c�
�.�����tӲ�������;���H"U� ��(V=���L���ml����t����G�Ut���|L����4�/*����"�t+9�5�L��K"k�k�j�+�_r��~�"�瀔1;6��Qe�ه�*��[S�?.�
>�|s�b�`�mK�m����t]h׽��"m�Z�xB�;�_0���]sw;?���w�u:<Vw,�r�b<��C��龇�R�c�����7?7nE�U�ac�F��X�����/U��c�ض��n������y��_� BhՑI��#�r�.���(�������pP��>_����$��:���*��4����P�
��Pdv��Q�-�L9`�co�\�)��~��1��3�Z �n&�"�m?[��HŃ�_�5(�O�D�y9JA�	)#�﯊4+�����9+��¹P;`<��a�z<<���em4}����g =�\�ߧ��U�ÏXU0{�V�BJ�*����*)I�|����������~��	=��,,C5H������l�;�M�l�����˔)̨o�Ш�����|j��H�'r����{ �B֩کe�҄e=Q�0y�o�.����!�n� ���bBF������S�&��f�|�ؒ�1��x�V��a�u�)pM�ֈ��\�0[����F;����g�Lw5���z�r�y�X�g�ֈd���Qy���9�HK]%^��`��
��9ޟ��kgѸۣ��(���\ ��f�i3߲�YU��à�p�N��q�%9hbm��ŝ(��tTݕ�J/ 9[P<���_��|��I^�R-g�%���q)h~����@�6��y3*3o%0]������;��	rr�6ȭ|�ُkh5vUC%�,���HU�h��F�����E-�Oӡ�3n���``,���
I^CNy���_��%���4P�����4�P��VZB$��^��3��$������e�sa�E�g<<7��Xc��z�f���ێ�H�Pm��=�2kx���9�\�K���w8�Lx����24 ��-aTվ�֟�ܰ���,�9˚���L����n�ḽۺe %�x�|�[�R��L<-����q�����&�Ĳ��m�9!������N�s6�T��C��Կ�c%�E�5~2��H#CyoY�(�xt`E��rI]d0{!�cP�v�H]-���뗬�"�w5|����u�=��l ���W�(ץ����򏎊ZY��BQt���qj~���L��Q�1D����=��E�&X�Y^�7�rF�����W�b 55
��G��OV���Dt��8׎��J���~y�����w6`�6c���� S�����L�H�/2�C��Q_�G�%p j�!q�q!:5n���u	"f:Z�T� �-Cܺ��������['�|%P98	di��CO�۫���/1XW� ��2^����TRo׏�~n!�W���+U����w�br�3�'WJΥA�q��:�46��F��% �D�v�.�;�`�U�	���G��)HriB/�1a+��^
+p�ڟ��:PDS���	���x'Tp���lNuX$��ou}��j>@���x	�R՜{�B�1!��y"�&�sY\F��}�L�I�4��P��!����6�$m���`/!��-��N�:dG?���8����4��R<x�<���	�L��2$ŷ�-�Qo��+9�����)��ē�װϻ��B�s�kǲ��M�e�-�\�f��uv�8T��	�ͤ�w���,����pr�Еة�=3�F��1]��.� �ꏲNƥX�N��5�w?
I<��;�.�S��u.��=��GAt�ݰ�^��]+�%IN� ˹����G�m�:�>�.	�;ګ	���w�g�^p*f	�ҥ)���JF�3�T0k ���m��Oi:Zd��Rl�n�>3qnB�~\�Y��~j���"�0���ˬ���6�����B ��/d�I�;o
Fwgi�^���u53�����7�������H��W��x��ߞ܍��|}"���^'�.}g���E3[���S
]�NHP���2lDeC�e"�.�K��f+Y� �$�=O�;Q!=��l�Ź=��f�8���[�C�&f�f7�Yy�K2�itP��q�Ztc�!dVw��i���fc�F�4R| 3�ѧ�c���-ML���ȡ��^�j�[�S;�,)�E���Q�e	6�6 5eX�>���=	�'�Z%6���Ҙ��_@|�c
�&SG���!t��D]W`!�YͭU��^�DL~�X��<��tr{[[�Wz�[O��j����\�߮�Kl��9��";ag.H�h�ِ��� ���;�S��V�����Kg���)܂esxr�(�*��ΜK���<���C�e�S�%8�o]�:����2w���Lm��
�i���w�5��Ś\���H�\s���L�^��<?��0$�$[�|�̫�91[�9Ul�������C%U)(��]Ӯx��aS�u�1����M���V8��l�D^��[�_��b�[$N�K�[3�:_Ed����d�"Y��;��� �
�Q� �]�����	i��O�?�z��5)�� 0�?4�&{1 M_:6���P1����Ve#��EfIM��ZE�ը��\�2��>rӱܥL9�	��,�q�'h���]���!H�gmG�?���RX1N�?�
2t���%(U����?z����l���j+�Ӟ����rԚ^$%�=�>Ia�/�R}�50��b�o-�|Uj��h�XlxVHYEB    fa00    14b0�H���4'��*�a�I�?z�c�W.#SO|����.vfmN�R`�n������W�0��Ӂ�ƒz-"P��45������k$�}2bҳ3��g�N�f���W!"� X;����(l�?f�_Q�: �g���~v+�i�ؙ/�4�W���2fY�`�_�zz_�F��7��߬�	&oΈ/7�W_�3����~B�_�|7��R	>�G�|��f��ӎ��s�f믡c<��,{�$g���~8��{`8VbE�u��Γ�$�J[�zܙ�n��Վ�.�߀y�b�8��~�������f����*��ry��u&��bl5���D�+�s�t�����/�s\�%SiH���5�������<EL�R����]���W�HV:3�ea�Ǌ?�	��MV��\���J��h���L8S {�=P���^�L����w��#)N��z$g] $؝���6g���]���F��m����O)^߽2���!�p^��̳��ӔJ��(oy�P�A���ح�GR�/���ǁh��s�`�w�e"]��r��x|�fK�Q�D���+*3ʣ0y��q�W<;���P�?�g��YZ�E���5�yq�bk+���Seu�㩐��|�?f���o"u5��QN���9'Ƽ������c<w�]I�]�Xi��'G��,0	�HnF&��*�`��%��q����� .R���2�L��`�/�=�Du+O��񿻱U�}ZZx�g�s��I�����X��g&{�.���9�B��=ŷ�����V;��H
�Q��H
[�v	.��ah����	��p�Z���A�[�}��D6L���
o�T�9�FA=�ZaK)q>���k�BI��O���]����B���*�YV�jU3�
���+m��{�b�[<$����ws�rƇ�J���y���[�"��57v�7��8�������ʣ��W���iA�΋�ħ�R��׃4�U`e{؛#Y��׍��l�GM^��0�m�S}�Y��$�Ղ��@BKZ��e�f������+P���fyٱx��i#�"e� ��Wr^�\l5�l7�B�w��k�"�M�ȟ6�T����%	`�X)ѻ�	����u��|��uy�TxsI_B�0�b�hZ&�����e�xF(��ˋÓ�:|���n��!@6�O���~)�<����.� V���6�{o,���J�ꩾ�=m�Fga<7��'�P@kV�#n?0�^B	���.��A�>R�'���3U�i��q���e�nr)fAh�ۘ���ܬ
	D7͖�Z�E�FJ)�v�V�����w��6P��Abɘ@��U	�*��'��)�����v�GC$Q��ME�'�7w��}R��=�����C�|Ŗ��7�%)7�k��A9)�+��^g��LAy���ϿH'�*\b�4��f��<�P�Qp�i��;�U�8>��,�u�=!*�o�}r���W�n)��#O���Mu�o�o:�t���=��z���M6딟9� ��#P:�?)eNә7^ ��G��`�+�HxF"���OSw�U�n���G<]��)�(e�8Mt+Ka�s��s�[�aH���r}�/'��x|[�,�������4�a\8`����Ε���qF���z�f�6�������b�ڎ�KesE�] w��~u�3z�N�v�&/¾3I�H#�|N����z��QZې�Dc�b�u��?1�qP�{e�i�~��;;M&R5�r��΄����6`�����A�]�q`s��Id�^�n]��u^��w5�����/�Y���0���au�7>0���&z/�`�4/�����Q�enjBa5ۂg`���"��RdBI(��SԐ��VLW�ق+3�{[�J�,Yv�|t#D'{g�!zF���Le�
�����F�i����Ԋ����M�ֈ:�,Q��, �E0Oq��҂�#�$7��-;��i�I��Գ�a�����0\N������i�N����y�eg�O,3�O� ����A� N5[}a�,؄�`e�9�h��
\���s2c��pѱۜH�V���\i?���/��r�G(
�.���TNňT?��t��ZV�J� �59��E&��|�!��� ��7��д�E�<��Nd-o��M�Z�o��,P�7�5�'�BJ��XÐZZ��F$oo�|0��\�����ţ'�7RɮX~��n#��)�M�ockƭ���z�3 ��#��G�!��$>������n�\��27L��NB[w�跷�Yw֬�,�3{�<ʽ��~���ʓe�m��%���Z���@��r?����2kNlk��H�O�Rv�xt#�������3/�Ӿ IU��g٢�1&[���E	���/�2\_g% 0�4\���D��j�+�9��-G�{��yu�tP*�E@��}���Ü�~�9�d��M��p^�����O��
��N�qO�g�$*���hb?�p�K���F��h�0?��$��hz*0)�����*�:J`WZ�{���5�i֙��&*$|��9�x�ۛ���I�x���,"���>zNP�5}�dM5�J(�e�!���R�����2ڃ�3�./�eG�ׁK�#���:{·=��v��}K�lb��m��>hn@��Եa�-X�	���(��R�ѩ���m�Ni�+:�\ޏ�8�D$�Z_�OU����V$-f���⢤Ʊ�Y�s�,�6\��s�xw�r3!3�HRB%LqWe�\�=�����cv����X���m�4�7�ю��޽^��U���/�����M���ո�}JӗfʶK��7���E2���f���]�	P�%�8�[��)�s�g��K� Q�y .ET;��l��z�p�ih�;y��
^X_O�<�:�</�e8��E�(&�a��Y��}	R��#K�8/=cJ���Q��P�Ѧ�^vn��M������"
��e;�F�+4(p�p�:����X�@\ϱ&�fp��PC5�'�!�V���w'��ݍ�R��1ള�i���p�ނy1;�kn��PV_�&� ��`�͗e9*ʀA�Bq�y�&5����9K	���,�(M��tn߸"���6�"�m�k�o���j'0.w��l��A���`�#�A�;3ĶR/1{f����
ϴ=ڣn�e�Q���j�w�p��|pf�*�1,�jw`e��v��.F�^������pc�S���S�C�f��L�����!�@CO�Ѧh�P@^v����>��`�X�#[n�;�y��R�BB��l̗�3�n%QCY�L��F�W�J�]s��ھ����Ǣ�O%��xI9�����:3!2�f�~���Q��h�K�#N��*��(���j�f��7b�H�="��ʯ������XЎ���e�hެ�^s��r+����A���R���(f��CD��RL��z1Xet%�Z�g.��eZ�������p����n�T3A��x-Y[�7��7�D9�2�4cm48�mJ������R��sQ�!�?N�}v�-33S�`���{�.��粐�~o�M�4MN�@;�h�E!ɹ<|l�l�=V�ŷɭ��wDXp0�yo�[9�c24G�?�4i�ՋU�u	׌�%[MԺG4��ed����
!�+l8�����.��/;�_�>�Z�Ɩ9_
-)-����(���V�$68 ��I��ܿ�N�0��
}����^T�/��(�` �A��B���w��
��5@���!��e�s�^&�ŪjKw�X۴�3'|
E�C���2�/���4A���B�:���|���OZB�`Uܝ,OI�K�=�^f\����`�#�bD��g�F�geXCs���E��	�\�l<��B��7�|d��n�k���s�A?iR<��`E�m\�?���`�9 �n��#�ߩlJU���?M��_����sf��MFSE��c���2m-�s���m2�JP3GF#��4v}ɇٍ
Ȥ2��Q�7���mᷢ�w���y<�L����+/Tƽ�A歒'Ï��	�s� r��>���Tgਜ਼��Dm��(�O(6+�!��c���f��O�$�UO�T*,ˑ�s䘙�ôr`DW���#^�
V�21p�{V)���yj;���|R~⡂Ǥ��k����[֕�v�sr���"Yvؗ��l:��\�༂x�]�����H�sm���8�p�(F1��Q������xM�i���x��|0T���i9�ͅ����j^�=��SD�Cc�F����Z𴟥�:;R�[�����"�)��"N��F�	}�ٲjH%��ė��~�!��$��$#B|>ߞ�%fi� ��1���0m$�>T/�mD|��d ��}�y�4G �?0	��lR`H���ȧu��<���9j�����m�Bz3��ɻ�$��`�w�nyI��y���kX�i�����I�[!���o)����I���2;����<;�����O�)�[�Э� ���=��<���y`k�����&%�]�"��Ƌ�y3��Q��*��Lz���#>>滌<��.�\?l������Oo�V�?���s��c\[�@n��ȴ9@��+��YKݪ����h������w���*�g������!���8[CC��4���9�_���
#�?B�2��Y�U��et�L�l�d+��?wWd����Y��i?Cr ����3�N3d����ob��l�o`w�|��u�Qr�n���O?/×%μ��I�ڋ2FԬ-o8	ZV`6]�6��v�F-.��C+���u�����J�n�,w�9�G�'�'	޾�Ҹ���1��=�0WH�ƕfy�A�f���R�F�C�Ȼ��0e<v��tArP ���ᅥ���Z���q��
�7����[�6A�mP��V �	.�b��8������?��()i�'uKAK�!�B��a���D^��������?��N6Kp��{��~$��"<�DRe�u�kR86\��5��Ӻ��O.C�T�,g���8���N�z�T�^��X�L>/>roe&8զ!.�L�P(\�/��6�L7�.O$"�z�6ĕ)#�� 0!F+��y�g���݋������sw�n��O/ie��od�Oj2�I�rt��5R��¢X��p�F��ą���nj�c�T���o����1���B�4E������<��LOW �EI(�<iќo��$1mI�MXlxVHYEB    fa00    1880a�oOr_���\8���;�!KO(�s���.@а���ӊ���R�`�Z��(�]T3��y�P�nң¾�8�2k;
�A��ڍ�`(��E[d1�O�"����r�;����/��a��g��H����������Ժ~�|:��>�������!)�o��S (=�A_�
|�+��-N��+{�?#/��5����7�Q���&��:pi�������ȏyj`���Jޞ�ꥃ�B���՜;(�; �좠k�
�UB*g�d���+8=�Q��Yђ{�;����Ua��;��x��0�#�鱗��7�˾ޓK�	rX�C:�u��g�u��r�M0�$�G#uJ����걟=�Z	dj�#��|�tg�
R�:�Gϛj�0l��4�������v �|'�9O�̅/�Z! Vn�&Ғ�j��_�����a~P�tՀ���\����iϮe��t:�&7 ��3����nS��n��_�D}s��\h�S��!����L�ojJ���)'�q)���M�$��A�#���)��xUos�c���2��["�O��O���1<�t���p�{�B&ۢ��Ѿt�y��4�a��k�eP.#ƨe�-�`�^�z7H�4�J���zW��6>�L��H=��zVcP�рRTx�����%��v�@J:d)��|�����id�G����IG�V��'���� ��7�8Z�:�����x�u]���c�!m�(?��"��������ueL`����Q;��ğo���X?�I�oB����p�NKA�8+\�@���	�(���E�ٺEd:�Ϧo�~%
���\E�k�m�ҷ��
<��cEĪC��N��7Y���䲀���\���}�n�C|ϱ�\��Ph�{K��#2r��σ�"g�P�M��B1�����.dn�D�|�^��ʽ�ļ����v��û)������������P�����{+8�tm+�W�A�A�{/�
tn�4V���pP��ƌ���Ϋ�F��8FɊ7���K=
�Vn{��S��f���qf�LB���p˔Q���{d��q�p�KXU��AQ>4����@���tv���WQ�0���pP�{�#���ܝ4v>�S`�45�O������;S��z��-���S��`g���-/���#}A�~2�]Z;>���3Kq��"R����I��Q�����qB�B@-�cp�>�#��%[L!Q@�E���+~�M?�a�J���|iU��PG#��cQ��	g�y�T�p�أ�4���o&��4�>�L�`4M� 
G;/]�^*jLY��.�4��k� �Ps�$�
"M[MK��ۤ��z8Ї���Ͼ��K_��c�tف�
�����,`S����/�+qik,����A"�G�������ku�h�h�-�3�<�iƍ�YZ��\9ž�Rt�=�``>I���ʤ��Vï����9�^�_��I��n��i�"@�th�FU��:���⏏
3zL;6'�Q� ��� ��Uf���`7D��& 3����V�����:$�H�H�I?��.�ߎ��#��43u��]�f��1�H��L�GC��#8F{>�]j`��/@�j��e��D^�J��n�c�hk������S$ٯ"�},�3�? ����Ҍb62��y�G�~�^��.0+!Ҫ�AC��/��������/���(D�h�Z�J��(�'�Q�	��yn˂3��q�K�`��~�i::�荚���@`��֌��an�ޯ���88�o����u&�!��l<�lw��ެ�����ߒn���H����	!��h�
�.�_%^Y��~�>����A�� NHP����_��AL�V��0���Rx%��=1��Q��������t}-:���}���62d�H�L�� ��/�H[��/�`B&%���\N�(��G?�?-=)c�q��F��2Ԉ�d��6������4�o��)W���j����W��uP���jhQ�[��V�QԺ;	
�f���C�esJK5QJ��	��T�}��9���9��"�U�6������� Q�[}�TG���q�%Y���h��뛳����0价c���9�d���>�o[ǝ*.ޠ�����p�:���lp �t����}걘tj�2��gU��
�U��D����� �GL+K˾���RȎ�#px���1���6`��ԡ~	��Wn �㱐D�:J�l</5��v+\�V�Qс�Oƙo���3�y�N�������Af�M�i%�����D�-?$%�t�u$�OْH��@U���Nky�� �V���������-�oӺ�q�^�ݪт�!�3���̐�������:F��s�c�}��`��
��D,_vέN����Z�Y{}f���Ȩ[�ß�3��N��_K;>S���ng�H���\V�>Y�yR=8���&�gB�U9���yy)Ջ�,Z8E���:�`�������p
�]�C7 ������g���:�䲈g1-���?��^��ok>����^`�[�Rz�-�,��4�%�������9��Jơ4p�L�ظ�e���!�
fع	n�8��j�i L�{�FQ���ц!;��]R��Z'���RS��.�|���K�Y��|$7���Ʃ$_������ ����17�-�Th�K�M�ǳC_��,Be�b���!2�|g�tm)�0q��?㫛p����Ż!|}ǆN�!�a�)־t9�co�`�0?k���o���UK���s�ݯ� �CT��JY��#~_t0̐�+MV$����ŶG�$5Ĭ��ǰ�T ���c��:�Ӈ@\Kg�@T@�ȱ����+�Y�o��K~��Zp�[+��/NY1H�6��j�����hn��#9�SFBI�@y��繘��.W��������geX��k�$V�(�XHE>�S�hq���1~���
t��S6��%�Σݛޒ�tڄ#�����g[��y��>JG��J��]� �l`����bX�w�0
���-cD̀�/���6蹓G����$reμ���\���v����J.����-���� �O���hS+�ݛ��kƉ)����ʎ�Cxh�:�a���@�����8{��l�.�>߆b ��m��&���Coq-|�3�`�[Nb��Ee�}$��{���se@f�q�Q)��4Ij�r:�:���O�V�
��=�(h�^H�Cu ��S���R,}L���jl����R�4"�P��*���꺫t�8z>�O��C��΢G�.envy�޷'���(Ȕ$���S����U�Q�˗q�z� ދT��je�n��#�����U�nɎ퍩�"M�&�6`��$�!�MFe�e������K¶9�geb/Z���@���aג��'{DgU�W@����R��'�%M���O��%�&9��Z��]�WKn��ָ�cGm�/��/���p�(�.^���xB���ދFv�O���k��4�hu5n����<}X���嚼�� Ɇ��S��l�Â��*V�y�c3)�X/c�Qa���CMY@����3�X(J	����(/z���*!JZ�B�[}�<��Q_e3�s��(�Ƶ\{M|H�� ���h�J���f�r˨|5l�= I�ה��mӔ������9��I�x��� ���\������`�tv8Ab��ي�a5Vh�[�WՈU>�mӐ�E�� � �+@~�O�[���yI����S5��TA����4q(�vB��I�>G�(�B���g^�X�Dh6]g������j	W46{���u����Mr,��^9����)�� ˽�)^p�Cj�e���	훏M��U��XJb�؛:t����D8ȿ��34�p��t�!RkYC�U�ل�K1��i�i�@���+D����H���(~K��|()Щ���5�h*�M⥁Ml�zh�aqʼC7n��n�59��L��2���'`��Z(y���b¥E���[��`�҂?oR�^�*j�p�b`�V�!��~��?��=h�f�����cm�Ԙ���"�<9�/�	n� �d��/}.�j��k�a)s�-,���bC�tz^mCl�1vE(<".��eS��~ ��>`i�l�GScdg�g��z���ZYu�ڱ+tvϪ^�4(���2x��mC�Y1����7����Z�c��Ȉ�,�:���,�3�8��H�Sz�:rJcƇ�W�&d�g��P�Ϗ~�RѳfÎ�#1�oN
��[2�{�r�\/��9a��	`�bq߀f�g�^������J���̝�[��䊨����?Av�WF�8R�Vu��Q]i�=��8%����g�~Q��fÇV���oM���5�8�cw,l^�y±0E������5ǉ#���"�M��E�sr5^yI��f�-er�����
�ub�HA���΀��_�
�����9!�%�Ӥ�.�ʱ�����JZ="%'`���ԕa@���cr��/}.�?/�;���_�5�e�1X�������Gޙ�_���8�榸(����r߳��ߏ�I�8��k��.F���� !�	:�Kq�m�7�&��z���w���Z�S��5N{TQdy�%�o��=>83�zA���H�d\�>�
��D�r�c��������������e�d;��5�wc$Ҷ���/.�<¿9.w����]0�{���O�VcU�bl��x�޿���rb��P�1Y	�{���������/��H�~*Om�$�t9�p�[ġ���|��9x�F�S��@�e�C�������5�V���]���Qv�V�tg%�x�����/"��),�)�]������/@�.�� _O�k �H����8z �$w�B,3|Xv:�q�; N����6�u�ă�6K=�毚s�`�؈U^�eq�LY(�*�N�����b�3����� ɮ�uF��,�Ek�N	}~��0,/������t��E+iG���w��C�����P	�˦Ϩ�m�+��9L��\T��P-�F7�??�@��(n1po`�+������T����,[y"@����J�������I&��%���
�.���H߶����}�����7�u�t�C;��� ��_�Ғ!B��5�vM�H<�p�?��� [�̫��U�U�����Z;��Ʀ�qۃ)6����F����C�#�Agt]X��Q-��4�ߋ�W�Ǎ.��/E%o�A���<FO���><V�S�8ڳ��qde�8�@��M��a"�
�š6�V;��f�9�?��C,�S�Qd�`��lO����ά"��8TX�4ΏKȈk-7���ԁ�-m��C(��;G\+��N�}��S�8�9�T�m���a6���{,ПS��֤>��#����&w�1�=
=��!��s�{���E�}&����V�_��!�$Mz�
����E�(���,ƴSw��t���>��4��?�[.���Y�ALV�l��sY�I�cZ}&t�����˵U�TR9�\�6�k�Ib^���%}QJ7-g�.��AZ2����ծ���]4�1��y��ڕ~�ۧ�u!��S�����yͦeV`�qM���{*_���ZM��Җv�qV;!e�0�z�����g�9È�A[_
�t倮��+��hg�y�sjF�B%w�0��Թ�ú��~�a�j���^�O΁ι	�Cps׫!����'�����pJ$�H��
�R	�C��uN�����P�E���C�1o5)��o��O�"E�eE���O'&S4[j�@��Z�e
�%�I�k�@9���fQ?���D׭�T:���?ME�����g�'n���oÂ�C[�`k�g�������"FO�>�5 �?o����	­�w�.M�:-�j�^���̦=�Vf/���&��>��s����
��Re��)WUQ��ˌb�cH�$B�P
ɗ\q]��2�)��W�@�ʐ�\y��k��Q�?J��N��a�o]���O�h1ԣd_���z�����0��)��ˀ��B��5����0㙮��/ܻ#���O�L�� O�r}./��EK�w�,�+υ`�F���i(�O^t����ǹ���ZH₳�L�/od�Gי�&��+-�h��>[�~*f�s�[t��R٦�-��1��9�{��ѻ]��$��L����H�b��[��Hj��yu2M&j�=�5XlxVHYEB    fa00    1910� ��QΈ7@>�	�xS�OL��N��b�
I G㳈�}�|*\b�|�H���2�~���:���]aR���O���#�@��-�x�tx��y�P�� �	#�z�յd�!2t���n
'��uH����;����W������ė�Yyn�����=d.��9>lN�WA-;��Ue+�����U�-�����|�:�{�}����W(��r�A���|e�m��;���<q��,�-��ﷺvP�$E_+��V
��?	#�D���2��cm0Oa�Ȼ����>�%=��^f�|jHY4*�Q_f�K!��QLco����˥G>�9?ɻՃ�IY ]h�����:��W����Zic���,a��Css�Ȯe�4�I�g��0�qw����6c�k�
��?�6���?,�V���VS�~�V�)H�R���� /�l�]��98�h�j,*�۰bXРh�5���K���đP��<|ҳ���AFQmP�>���>�-a�C�-��YD��hf�0�sG>�+�O��ݦ����X��.�<��H/�,�P��HLӁ�@�l���~u��=�������� �\��vǱ(C�D���{�z+�#�2��R��&�'�%��6?Hy�u�,f��7���ük��qhWgO!,t^)�M(��RI/��E�r"ϟص'a3K�p���~�׍b-���-ս�x�� ��� �B�¯�ý�D逹��Í�l�}���5���b$^�QFIxx	�L9��B-�Ǎ�\EV�����
T��uǪY<�`p-�ki�����z��n��K����n|1븃5�`��.Kǫ�8#ҟʤ�C��h>�h��z�߸��<�9X�b�͗	ѷu�J��D���c�aۜ�����#A�ن��*^�tٔ�
L��ig@��w*�;Z���9��W��p`�.��Tv��h�E*�$4	xr!��6����YImc�v�ͲN��DT�<İlFb%�كo$'K����V�+GE�[�J��YL�Jң�%�,��Q:9	�!�Ox�?#B�^#�k]�|�Bmpi�;���D�J��U��\|MdF�U�+�u܂��4�~iL�g`v\c��S+n��}�8�`hf��<Y	UeeJ	���2Oԃ����Ԉ[c��c4=}�Bo]�nA���Ri]Y�kÒༀ��H��z��_#�9?v:��V�,Y��lZMxn�kX!3W�4'�DK��Q�R���-&[ ��f�WG��_�7qE�{o�\�Fl�K$\������Rm�,���� 1��o��i�µ�B<�ŵ��+q~{O�=;#�C{�<QU�\�1ܱn��zѤ��Y��8�^xB�q-?-ϞR�~�7'�l 鵹�/B��7�K3%���%/�K�Lg8�X �gl����b����BjB��xV��A�O�i���/�e�U`�!�ZTk���Y��#kn `��A$|�`�������<v���ӽ�A5���D�h��s2\JRx냝��!]ahC��G���εH�>���UǕ;�$h�
Q� 5oTK��|���O��� r��|l@�(�u�",\P�91�j1g*�!�\���^N_7D-0�lC@��dŁ�16��
9nW�G|��F94�9�n�H��F���ޖ��,��J%�7��y���pA��%��!�>��/,��q2@�oP�t"���3O����{�w��.8\퀚EBF(��O}��<��7�=Kq�;��d���l�~��I�v�V;%�W��@��F����K�u��f�~���i�S3�s^g.M���x���߅���#yV�8.���8�=���ʦ%Lܱ�%#D���B��$�y�b)�O��~䔗5ʽ#�g)�>���9/)Ez�r�dcI��$�y �$�̓��r?t��uKn�w��+��s\d��S�bM��9�3�b֪U�r)t6g�3� HY"gdR
�@�E5`�����Կ�����Y�̃�jP% �*l������P�C������q<a1�(W���uz�F$�g���N�N���ӕ�Y�J��l*hh;��pvx8ӝ���Ѭ����b�`��N���@�!'?'u��c�l�=@m_n}��aK�ڊ_mI��]���H���.�C�{�
7י4��V�b���T�����g憻���|���3�נ"[�P�M,#������Y���I#��C�f�Y�Qd�I�'�����[~��u��S8X�9=!��jUq�����{#@�A��I�B$�RhA�w���=�؝�<HaKI�(w����Zv��3��œ�a����esB�bd�ƈ�e�/���ۙ�������S-#�^��t������0�����>�䝯z�M\�r	Z�k��ܭ�I�ҿETn*�%87����R��z-TWrR�.�raԸ[��-��*������M��X���r۱������a�h�R��K�d�	��`�>�u|�*�"p�T� ��z���0U3и%�G�F8�3S�e�Ow�^H_��Vhиs�u��pFC�r�m�C'L��r���)j���Y4�!ԡ[�:� �������|�[�*m�^��e�a�����������JG��3�D�x(�lE漱0WV�II
i��!���-��f�k� '�҅�&���z�q�ik���_����UgbJV␐	��Y���c�a�����e�2�_�k��ڷ�fP�Y�zU���0�w�� �W����	���-��ߣ�.N �3hXA7�c�:��	=Q�-E�DI�M]�¬|�T��/h}�bP��)��k���a����H^���u-s���
�?�)�v���J��Ghc�mX3
�)Q/B�ș{�ER���R��Ǩ���J�,>�G�(����m<i\ EL<\��-ok��t���� ;[]33z��F����_�$v�zo���P�,9�V��fzt���k�cږ�`�F�y U�1�/��.*�3�dX������ؑ����,:���r[K�����'$�����f�BKU��%N����~�㐸�Z���Ne��J�݌�f�|�Rs
[W�9{����z���L�m�p�c۬�8�[����eH�+����dZ_����R(V���S8��܈�� iw�(��oa!§� ?%�N���ƃ�&�4�5�4�&o��8���'�b̤7���9�fT���a��������B�Gq�(,�q�(M1E�E/u�~��� �����g/eºnHE�&b8�C��-�����"Mf	%�4se��tզ����J�p!����8]����Н�I�OO���Ác%iF�Ӟ���HB�+��"� �X�shf]�a��_�m%�G�@
]+�$"B����N*���Њ���N,�K?~ݚA��,q(�>��q���A�O�qę�f�9��߆Z-Y���Sq10�x��ل�W��e�ڸ�����R�����F���O�	��@&gv6OF ��l(q��j}U ѭ��󆺈�b��=a�/x�^AtXU�|�u�w'�*�Of�T���}�'ڂ�z�r�!�ïh�U�=�7�mx����\@C��k�R���c��� ^te:8�3���m��i��k��Iۉ��o�9�ٟ�ˈ�� ��4���[�Ԅk�'����N��F!�5�]ƩS*��k�7��j��ӧ�B�q��t�V�Y���Bw��e7��i��:�!|�_r�	��
���x��é����ٌc���B�K�����fƚSֶ����{���K���%a�%6�][���:$5Xm�ɴ0m��N�U���m-�)D ~/�b\P2�<_胥����y��`�c_j�/��ύ/�Ѩ�.���B�<��=k
�t���Ҙt^��<�Dɠ�Ƶ�K	5a�|���cQ`�	N��7>V$d��9�[���h4@F��q;��0�S�80��bn��o#M�3"N�o��Y9Y�<�B"��r�U�<�/���O��gDE�x�y�u_�C���9�2�����0p\��ᦷ��骪q�����(���H��P�E����p#�s�P��.�W��k�K��@�/�0w����uQqW��ƩՅo�ӣ}�f3!�,ÿ.��yQ��^�u�|��+0���Ə�O�d�l�B�:�r��g�?*�Y����?Dp��F�y>d)�v�Qd�cX�÷,��Y�{�5h/��@<�����F�)5?
V��=��b 2���~wr`dȗx���7���Ւ^�{�y�^��ɩ^��}�;$ᦳ�V;Y�j�z-�/��КG<	�(Zr�2�J��C������J�I�i�����\92��HeA�=R]m~��_�k˛$(׶�d*�r��e.�3ݻp�~ф_�tW}PZ���%/3<��R��L��H�u�LM��Y�SW�3&��X�	e�-za`��?���{���ZR$�"7�$�I�[H�zo �CӚ�8C�Á`�M\�$<�����e��&ˢG���&mp�� �1b<��V'���Xm2L>u�:5H$������l�t�de��ʡ����*zj�N`���F�Y��;3i��p���h�2˃���Y��⿔faX7ƛ����+�Z������>�u%x�X(r���ԏ�����d��³��NW�z|�S��l��j!�����G�����!�i7هM��a��F���:��#��KM���kf�B�+���9󘅄>e$Q��/�r�rn> X��l!emG�<�k�t4�yޏ�
�����<֕�����K6���i?<<���:��_���LZ�hS
�h��d'+�(@��!� ��� ��b�R����Rm�c�S�'�D=��c$ƀE%zk��zG�c�O��o	��� :ak�5����,���5ƀ���/(No2�d?}x�-E��L~ ���οsjM��A�7��*�?�ܼ\e،}��7�}]�A�0��1Z��g��n���[�i�5N36�r_���5ԯ>Ι�sk��{��vW@m���}6*� �]�L7��K���a���T;R��Qu���]��)�N f�@ ��A�0 EA�Qe��blҢ!N?����klh�<o*r�vp��`{�#*�gF�H8�k[�K�v6�l]���X=�.��Gg!/�>�Ns|9=� =SDy�<N�δ¯����g$��q'��|�䍻�f�aO�����ez��;���}K>Y
7�	m��J�.��v�<4`1�n#�f�*/G@0���'. <>�%���JM�=��'uRC��K�t��� _��1�A���xu�ڡ�������*��fΛ�%�ivŰ�pfQ����j���10{(k{�<�5�f�����gz�45�ОS�sa��Ӄ�6�r���p�|fT'��?���E����"��7���Yy��o��lM줹{5�=B��H<���"��7T"?����jxg�@�jo��w�?;=��B�@��N':�YBk��n��lf ۽[�]߯�X�d�(�K"�N>�͌it.S��ga�b����%�ޒ�E��9��<��MΪ��6h&�jd��l�1��KU���ۻB��3z�Qh���s�������m���� ��������wXP%�6���_��{i�(v���~`�*�Xw,L�ֵAw-+}�h=���j˙r@�#��|<��<��̒�C�wנ����/��ؤE�5�I���e!R���k�U* N�N�/��$�ɛ4eӳ��1��a*)�	�鮦�%C7w<��l;*�>�e�1RH�4�,�&��M���ۏ�JTi�K֬*�ʒ��8���;g��d���x
�	�%�-�yX� ^|������D��077h�N��Vb���n���T»L�YWdQ�'��CfaVe��V�@�s�qzu��*w4;�'�6s�^�y���m�Oq�ryڹ�	���y�wL�)i-�?Ǖ�]�~��=`�p���51���������؏kK�&Om�;Rj�i���pb�~;l@��P�\`�1��e��VD��ǂ���z�^���վ3���
$W�w�y�{���&�P�@�GZ�4�����BK��ϙ����竻�5��_�;��ƨ�����E2s�9@�va�����*to�Sx�N�����`��hDb�h#!�=}�S�n�؜��*!�P5�j���q��W� ����2d�n�K	���c$\i��ǥ��(%6�
���y��[�o��W��T�f�?�9�ي!�e��F����j2�$����N��J5A툥ʃ�S �S=έz�(�����Yx�
��q_T�8��q4ՆT�g�0��i.b휪V�|+^�m����L�w	�u�;+�4�I6��%XlxVHYEB    fa00    10e0Mdyk�WT�c9-R�uq0�Q8�B5:�Mw"��lx,rGz��/�)K�@ ��5�K�z�g�61����P�@�SKylH��_az��k&5�t��XX��Zr��{\xs~������~)�g�_��S1tn�π������\dC����d�li��B��@?� ��N�WuM��n�_?B�M�*z�/5k�c� ���Y�z�ֶT�Lis�
"$s�[Dް����;wu��Ł dc5���x�A��8�.Z���/��<~�[j�n�I���m-|�7u���F�ۉ���L���"U:@�p���<����!��-�U[�,"����I+������Ϗ_Ͻ�e�Ovl��2�L��.yG���o/�2.��i9#����̭Qqn]�8} y�4�#'�b\�s���0�N��JH����`�5W�-Q��E�h������$��5M$�����4^}B��c��<S��6�}��.l�?���ܚ�5*�A�R�H��%I#�j]ʔ�T�cL�?
�~k�\���Z�mtүx���`���|BJkQ�2����}5��H�*��τ�YA��D��%�b��dJaˌ�g�
_^�z6���k����23��t�p|�i�"�W]"��	��{hĽ��7Az��������b�Ò�˺⤣RP�
�őxC�c^�=� m���K�~�I��dy��%$������5�$�o��;jO/[�@E�7*M�A�i&Y{�|�T�n�h�u_`�^�"��]�S��f~���3D��7��J��NI�ˬA']�4ʐR�W�(���7ȕΆ|�X��>�-$���s�ĝ]?\1�����w3��{ܔ*i���y���x��'��C�z1]�e�j'a`���eE����qE�#t3D"^Nh�q5&2}�b�,t�W��y	~����2�/!u��'P�tz���WYs^P\j�o���-�\�2\��O&^k�mL�-P���Ϋ�����_T}�()P�}|�!m��۱���� �9fz��+��%4���Z��v��c&�޵�E�4��j��VE��&k����$�W�& �.��O+_23��>"Ј
2/Q	��N��V�U����4��*�f� �S�b�
ؿQ���?�q�����'?�9�.F���;)@��~�'�O�[�{aQ��мބ/Fb�kP��a��]&�b�3��hX	�0��Y��pv�!Du���ؾg
������\�[���MH^�q�5�l��5��Ja��Z��27�39J��-���˓�ӥ�͸,h/�b����������=c@V���	A���ƙ"zL~�?*`��R�#�$��%m�p�V��ye�^+��U�c����U��6��}uJ6~\��NYsO���Z�nܙ`Q`����^H����J���f$K�O�IW��?螡K:l�h	*ݿe��]�fmm�s�-�+Y�B��,a"���EK��B��w���Z����e���'@z�7�)�"�������J�2%s��P�A(���Ј�����3gg&�ߘ��Y�ou�)8��C5ҝ�k/;�uTdF�� �M	�Cȣ
��X��]	a����u���oSlŧ<��mn���t�M�?���6wX�f)u
yu�	)�D%�=��"��ωȺ�:�6?�Fݝ$]�c�W�dm{zC�}�ocG��{�(�Ҫy|�{a��v��/�c^ߔ"<؄�f=��_1�,"v=h����;D�I ?�ɚb�����>�
��vf��������`�K����q<�0��8�ao�f� 1�7TA
���Z^F/�����0T�0�[%�]�;*�
���'S{����˭�ۄ+�Lg�Xl�����:
��=�\i���z���{����;�Tϝ]CeM�39���k$����I1j���nu��X�m�Z0.��FKU����Hہ�������*�����k�k~�ȴ��3��Dљƭ�~�:*~��=8w͐�͞��j:6t6%�@$�Ր����P��H0� �`Kf�xKT~N�Lzp�;����a�1�b�4H*�����&�h��`rp�}���H�2�����_�������� �O��#��qڳHHfE�ם~�~u�6j25ʒ� �x2�IU7X��n+���q��	�(��Bx��<|o�	v�*
R�-%�{#��þ�萾J���0A��K���燠1����$jcowʓ��d�i�A��̃v]��ڱc]�~a��+�"Q�.Ժ�5qd�Md1���>�jᰛ$b݌{)�������r�Z"F�m�s/F�]�i�3�7���"̡�]!���C��>���(�UN��;*�U����%��nP���T8
�%5z���{`�v2��``���ް}:�8��#��@�H�=eH�c�c�O%�2������-D�$�.�̔�]Y����[U#���kC�e|&d��(�h&γ�$�pd�s��]�{!�p:�SBD������!B/`�g�H�̄��0g�ډ� �hE��d�:�C)�(��9���2��A_.�ф���$�	���q)��2�}[|��3����"n��u��S|�y��1u��M�-�^�m@Q�1 �i0s����\�f#�E�|m�t��8�.���vj�)Kj�zx�޴r��K��8V����/u�y 6��jz���	���p��z�2HeOEF����9s[g6�֮"j�3���*�eM��z�u�]��3d;Lqj�mI<ր�G����ԟmf�A�
�c}iß;�,>`��"�8��5N���Bb;�H�I�/�'dK[�?B8�Ac`�(��1~+�����P!�Je���NW�(t�J"��N����-p>����켱��*T#���o���HfV���H�Ɓյ���Ԝ(K+�F��t����J�i3��7t�v/Sl��\��t5��V���N�R�Ěa��^�aA���H���$Nbr�>_�	�{%<����* ��p�>R!GU�$����P��L����?~����~$�+�V$�3?���yNVg}G�&�kf2�p�綝�t�M��7�-�"Ĺ%=�>9������׼�@��+{@�v�+�Ht��l��Z%*:M�uT]t$����L9�����\��p���T���?���K��+����fۿ.o�m�\�r��!��ɕ&Lz�o��;�������Y~�W"A�=����+9��C:�ʖ�Kէ��>?��_�
�&"�ga�ρ�e+�3
.�1��0u�0s&�LM1��FN#က�j+!���~���Ͷg����݈�r��|���E7�'���^��f��S�ecf���mG�a��."���$Y� ,De/G8=#��Ɔ��/�~W� -a�C�N�:-�ķ�G�t^,3��f��-B�O�{ x�(?}E�t�1X섵�v!������=��8���x��O>���gG��p�@�,��K�(�p���
��Bt�J�����2>�Y��[����H���9e	��r���M��˃K3>m�j�A�,q�{�c����]�CTev���"|h�T(~���,ky3,��T�p���O���yr��u4�کđɵ2���8��daV�.W�uBE� s4_�L\:�3�W����L�ԙ ��y�3��H�?�.6uU�wЍ29���j����M%��C�ni�ĭ��7�]f��.��ͩS��L�����&��]�~���A��m����Jh'1#���5�\��yZ�`���v3�sv'�_j�Tv���/}ΈK4S���ڿ�-^��l��"�ݜB�/݊���,�3?�ɼ7�W7�ћ��{�=�h��'�؉�1w�7��>��3i�EWw���ν�z������;X��pd�,�2�� ��^(��j1���g�L0�A2Of�wx|C�� �;(e�� ��6H���m�r,L�lN!�;(����v�`�l���ĕ�zԆ�rl-�.�.�}
�c <�S�%9+n׷=h����RPоk�Kh)�89�S�"��[׷sd�9��b�=�*X����W,��+%R���\<��o��AS���eŴ�>=��@HJ'4��#�kji�����kQlP7�T�2F�r?N�(���E�J@���b��[}F`فc㕜��[�ks+���ᆩ:��O"��%�r^�U,p��f���^�rHp�X!�
چ �qb2�5*��vQ :��(�~�	џ�o��J���x�M��U�g'����
����ّ	+�,ީ?L�./ϕwc���PXlxVHYEB    fa00    1860Z���9�2�@S��W<�Ԋ��M3�>co��q;����^����9�����j-�ߥ��W!XUs�*L;�1�$�Vb����(>��9� '�!QI\�l[��
�w�����w���s�9%>��o���Y����ByT�I��G�uFK�L<o� ��#��w�[W�!�m8�8A/��x�.���%��
h��89������Dl�V�uM瞲+��35M+�2ק����dp	B���Y<S��(=�r�v`P,K��<��������V�y���.0[.I�lX���o�D��#��j˯(���Y�9�Un�%o�9����7Zo��޴���+$t��1_�]�p �qX4k��[�G{[I=��L���(]��kѩ̀G��j=�4��g�!�e6wY�t[aV=L��l�&..8�P������ID2�����K7(n`@���"�N�}sg}����x�R��f�~,�v��Q����;��<YL���˄v�L�c|Km�$�t;�=���=з�z{f7ǋm�l��z��R�h����g&l	�dac�`�l�]� ��+T�coD��\��y[X
.�����1:IryԏP��%���`
�<S�'n�՝Orx�r3U�N��J���08C���Q�8��]��W.�l #.H� \qe��Y���.�R�!}�5E��B���C��A�:/�c���&�؟�ۊMH�G�Z����hQ����5��b�a��,�I��B*�-�Z5?�$���ea�x@���^�cV�lb���ք��qYÈC����\�w���-	�!6� ��H�ō}p��ts������2��O����on�D�k��N�+�njT��ꥑ��e�^������[L�Q�8�Ӣ��++�_&R;��c���<�ؾ�ּP`�Ď�o=�_��jemUoLAr���`R3q,�a��X���2Vx>����JA�:���*�5����[��5�GϰI&8˳T
r�Enu�ٵ���;��-���O���ծ7�^'�'mP}J��(uF��1�:�C*5�8��O�
& eр1��%����QVi��`���`���t�4�BbQtxlߋ�pߛۇ�WG��X�R��݆o���U�:T��� ���r�.&�Ȧ[b���͞��EhH��D�bI}�y�����Jw�@�9��Q�7(��w��S���ڠ�0s��\�7�ٛ��B��rz�̉�Bj��L�a	�D�[OSH��Q�x@?R���f��:[1��M[doL+:��S����f��`�Gx::#��^��-U~ȵ��Pek�Bh�zI���Ef��<\��k�ĭOX��l�/0bۇ��Ѓ!v}~m)YG�a<`�c��<��	3�i#/�g���� ��cx=����U���a�=g��>���H!(P�]]�7�ЮC4����h�do/�>Y;���c7��:��L��*ԩ�_��P�VH���og���_TT�9���"���1�fE��P��������"�Bvtv.*.���4n�!R��2 'b�	;�.q�����j�
W壅(	1�����4�n�U�`:	�_!c ��/�@Vy��R7����1��S�	���1����'�h�Yj��rT�,eқ|i�ĝa����*R4�A�	2��8���讧��N��NN� ^�����ǴO+m߽��8#��v�6k�U�Y�	��V���38�P��P!9��A�!ͣg{�߈��j}�C�[��N��!����1@�ݘ0�:�o/�Rн��]{t��t���v�ӟ>�>�Ez���^����h�/T��lwl�]䋵q�|�eC�O�������h�x�Oo}���H��Sy�!m�ap5���C)|��4�2�Xy��l�ʍŢ�HI{�� /yry/g�ɔ5n3���/��=��"��	>����3��V~ۖ���F�H�	VV��(�������ڿՓ�}���Z��*�Ԏ�p�3>\6���(0H�cQ3�6�V�k}Ѫ�\�)��Vx��5����mV�3Y�Qjk�94ѭ@�ޓ-��.gD��<4K����i4��Y��6���h��^,�GʃP�}���СphDk��Z:�m�����|�_�!6��L�oY"�ɂ��%R3�矚Q�r��h�!I<̪)r&iDa��=u*���]4����!ɘ�}>^�3.�ܾeL���,���f��@�������!I^���g��g'�3P�)��X)�9�摩�{�
���d���n��S��Ϛmɾ�-=qѷ)||+�7�h�$6������U��#����-,�Z�=�f�Z6�����(��穈�
���D4�F1��R
umD�قBm^��E�3�݄3�{w[�o�F�.jD�,a�<֛(��Sȷp��Â-�i��'s��t���0���Z�az]�8��	D���]�D�pe�h��F�Du>G��qY��}�������3PoSa�Qf�ڬU��1)&��{	Q�ݗ=2]�ڞ2�{�.(��]3
K�����Ͳ����.Ƌ�% /ܟʒ��U�'inu��H�V&V�۪��	i'ө\e�������0|��$~��O��������ѷ�xw�tw	�~�
'@��B��s�s�@�49�a��Myń�Z+�fC�ju���{�Z��g�B�3�/��sM%�ґ�0UZ�0#�\\��l��3��q���	.@"�
�b֧)h�
q�ڸ��T�7�����
�L�(�YP3��@��8���*���ޏ^���"n�A�z������փ��z��R��(�����Dt��#ݽ�"ji��A���9�jD��J��< ��zy�����	�Ev�*�]G&U �Ƣ�����;���W����EdDAMDG����N��i�8�8�c�2*?k䟁W/��8��JQ�p7��k��eT��'{͢��N/đ�iI�ǚFaÞ\]Nt����z	���bi* �s�|�y��ȯr`��Yhp׬z�.n��W�z�l� gڱBu�[lJH\��ma��e��كN!4\z"��L�q?7P��2���K�J _ٙ�D u��ϓO��}�ź��w�φ�ǒ�l_�S��]9FX������Q#Saʝ�߽��#9�Y�GK��йu�cM�f˿Ap3)��hh��"ʚJ򺞼�����n7�aF��J?��ֽW5��?_��Ԁdu�F=bFHFlo��`EР;���]��H�A�H!�Ui��G��6��=�M�������jxާct�Q�e27S.(���.d�F��nY~�p�� �ɹ���c�$��$��%����[T�J��!�9}�!���� �=ג*�'" b�EP��nƕ��I/k������Kz�'�;�Ü�c�W[�Z�r��_��)�[�*>rN���d��e� ���	�=?�:��7�_�22���{iV�!ō�G�TOa���d=�t������r}ri��FSg�:��p���@u�^q�W^5�c�S�C�ꢕ�����6��������I��b�ű�~&�}2$7k�a"D�5w< '#�M��d���U\�0��- X�!Z��h�<b�c���O�.2�U^�ܨd<����y�[��K���Md%%�X�����#e�����H_u���u�Yt�PʖH`��ᙂ�p@5��Bt�~��3j����sl��s?7�D��a��P n/��m>d���p��A��8h=�?1-*���t����E�R6��d'|;�_y��5[���W�#��p�IG}4����، �l��H�X�j4o��`$��=J�&M=��`�i+��%l7�<��KX�=�,M�SK����,�M��o��gK����n�옹� �ݻ/}�Jġ�A��+Љ;h�YCDm�*�p�=D6����w��d���w���ĸ������{9G����Bo��Ì��պ�֘m1S;������_��	���V���};=ӣۺ�����.	�,3����5�V;� 3��2�!�!��0�c�mm��j�Z�`���#g��"ƃ�~t�=nx`]AW�B�BdtM5���3f0iU��TT�G����H��2K;����,�G���@c�2r�������;˼�
F�|�dH_V��X�0�\#(���=j�V�$�v�/�y��.j��N�'�<�	J��~��O`��C;�~iu,+���h�����1������&�T��-b���8g)����P�a���""?���
輎8�����)�+{������E�.�z ����2G%\5x'�J��Y����W�o��:M�L�W�<��[���~�h�2p�����l,���M>�o����Ƹ�gQ���%�xл ��{q���k��N��ۖ�	��k9αw��;0�:��_鑎yx?��H�1�*f��h�̸AUp������cR �%1ۄ��H�^N]����z��h�p��+�<3�E\g
�Rd拱	C���򾺘U�:b>Kf6w>w�A�~l���]]Ӵ}P7�^*ǥ\B�^����� l���J�%�̞��И@(�Lq�ܴ�o�����<s�4n4�(EP�����1����*��B��c,CߚYL�F��������xw7(
Oqu���e��4�*�	j�B=}��ތþ�<��L2���� �T�Ry0?ڣ#	Ȣ��f .�����	A�c��!LW�����%�d�'�K��0�����r��#
�y�R$ؖ��U��dT�{��?����*g�5��%8�N:�U�!��[��h��ϗ���o��%����,|N<W����77��d���Y��7��w�ƔCX\�%Ж���ܙ�@�0��M�]�����S.���\o!n�[�`�^,4|g�C�J�FnX�9���a��(�d/k�ȸ��i���2ı{��&zV��a��@�����W��3^�I<�����xɢ���M���>���f�JVT{�w��/���
���4���h�2�=;�V���V���9������V!��C�H�j¶�8����Gl��g�����&��4˶�Pb�9h'A!�ʂ�z\9����0�W��"C^n_�wD�dt��C�X
E���{��ArɊI�+���S��d�y�2!�T�]�K8T��ɠ���S���1�Zh�w�<9CS4L{���ź.�p�6%�*�̒:S�B�� �cO¶�R����*��N�[�!���j�^�h�A�j��a��A����,��M�#C�V	���y���yf��א�nTw��s[.�!��n�hgٰg���h.2
6�¯I���J5] $�8���\a�����ݰ��M�>;�����,��P�嚠�|�Js�|�6�So�fݽ�����=KF��2F�;���2��֠)Wv���� ���9Z�����j2��^i	aP-*�qd��r�k��;X�.��h�53������B9K����rDH�5��L4K��T!�*�ţ5,D�[�O����:�38:y���p>|�/=�:-$Ӳ)D�;9
V�%��Qg]&=O[�5l5Έ����tP�7g�7�;7ⷻ�5�Q���Y�мF�V"I_��gqb�=Xa!`˺U �qq��F�����A#s�KB\jf�dmW��'�o˼vq�$�����m2�{ƵW=테,P��`����S��2�P#�n�*q�l�f��6��v���Jtf���&��O��|�]Q1�dpq�<���C.}�~$���ǟQʨ����$��T���=�{D�8�Ţ���:�{�70ҧ��Scx��e���o���zk۠���t��@�-������γ?�,���x�o'���)�^��*'
�QX*qО=����H�ڝhC�]|ml`������ܘl�=1�&��*��t-n������g�tu�wĳ���7w6R\��0�߀g�>L��G>���ߔ��ӈ�J��O��w=�LB.��IV�I�my��O�^ܴ�'RP���>S���*^EIs��:	����4?cݥ?���ųtus��Y�Kr�	���"�҅{�I\�U��'�A_���[v�y��X��w��;�i��C̜cć�S7�
�M�=����g��fŜ
��S����Ii��"�)}׊�t�� ���YXlxVHYEB    fa00    1720媋`�������M'5����z#��7ݣĖ9D��\c6�V�+���?�{�w�9�S��[t�Sn�_f"�M(��0�W[��o�N��$�:���h�D�ȟU�s���C+Ah	Ȇ܂0���t����~H-wٷl�P	o$ެ��Z�t_��O_�]q�����;����	_q�/�aH�`:V���X�'�Se<W[�;������gY����(�k@�o:����J8;
vOp��
l���?�3���U����x&��vkP�`H@����E7g��Ē3�i�_��Š̬(\�TH~_[��n���>k���%��3 6� !L�ѐ�?��E�-�=�4d��;cZ�g��؅3˼Q9a[2m��>�ݥ�m��+R��qc���5l<�u��⇢�bI��X=p���w�X���ɟ��&߼Vq�߳ѳ�rI��~�kZ�^J��k�!���T�Id�fnK�u�>T>$��lxn�����\%j���6�&�\���ڵ�.r��zj��������Ku׼Jl��F|�@mF�`���*�O'jPĒe�X�=�lY�3�#�W��"߱�|�����=�Q@aDbS�j&I~fS�I	) ?"ᵸ���`�5�������~#8-�L����}��'�r��,f)8.�����94��$1��RL�%��y���Ut95��zo��d�Ҩ��˙���'�K6��}�o�-4��E�3�]��C���#d^��^ĕ����YT��}u뺧p�9Za�e�*I�\�mJT�s&zLO��������"l����L�15��uPQ�Y�HQ��,`����DU��cTA�
@h�����L�~���Ѱ�r���(��K�^�f^�,�
6�pG�G��c��
�S�)%	u��8�'Oa�"�b����Өu���:�������D:�m�(o���:�>V��'8�}NH:�Ƭ�������%���GB��݀6�U8�gq؜�I\d��#���]gC<m2������9���i���h�.)���1ɍ�`�w
�|<R���G��!��ȵF���hF,�E�σg	l"'����k�42�D�k�zl�M���#vJ�v��`���>C��:�1(��ǹ���"z
a%d�����&�n��%��UKéjdS�!�`[e�/�����WIX��}���r��G���G9���b
�ni] `�����`8r���zs	�	i�nX[Ӟ8����N3| ��&�	
�K�����.�ˡ���蝱�lx��~Z(�>N��u"�����Q�@\&M�h�"�'�43���dM����%����LӒ��r���M�t
6��N 6!Vyax�yc�wW��*�b��T�63E险��a�"7��.��2*�6�n3�?����z��
�_�b:���ko�5m�"��r�j1u����#�;E�%Xڱ7?=Ӎ4Zn��I]FR=j=2�1����4����p? ���=4O�a�����&hݮm��R�<����� �:�ഷ����V�J�����{::o���~��?�I�<p�Ę"aCZ�(����\� ����&�f�\F1G��siwܽF�3�Y�c\^%V&��E�f' �
�n���K���'^Ĺ���7�_Е�/ħgI0����'?�������$����驓$;��~�-��ٞ����]�sn��Bj�����!Q���7WK���+�0���4�-զ�Ը����N��P��򌞦��G�Z7��f
V�=,��d��}�U��S��*=}���jI���f�&������oi;EU����a`����Vl���VO���Bp9�c-9�hr��Rt��'�0*���+K�O�M���oկ�;�NC�by7�"a��U�����L�*�[5e�8�]��^�F#.��:p-������U�5�������4���#Г�Bad��>1��9��ۏ�4�J��ر ����k�RU ��"��J�=ա0$!���;S�+O�A1�rb�"˯r9J�?�Y�1:fN�sU�zYSM�p���+F���������Z��Z>ᖙHa���x��ՃR���.b$~��;Oe�)�A��c�c�3�ta����q�º�c�<9���<ie�C�A~7/�K���4���샅6��h�`x���m�J@N���cS0�U\`t���u�c�����sy��l�܀�h��r����U�=�۹�E�["��ˠ�a=Ӥ�l �4�F<��|��Ev���8�P�"U
E�+ܕl�bV�$U��T�2{C�[�i��T�ո�7����g�/l$Y7!#E�m$�Q��݊�R���S�ae��G�ߪBk�6�,��?�H��݁��N�u8�I�ʸ^�ڸ�oh[!�9�����Y�R����*{seG��R�mT��s�K���7;P��/n�����F9���I�����"���Q��8.I�������[���^u^��ۅ�)�Fא����a"�Ev:���қ�t�x���]�)/$��>��@����C����o:�L��z���X���ꎼ�!x�8�0w�s�>&2��3�q=�-��F>ݸDO��,�b�p@��N�U�Cb0��z+��B� *.����j��ەt:�=�!��g���7�h�xQ+��P��@m���Qd�#�l��)�`C��2.�?�
qK���1�Q�[� bŐ��œ�rH�&�[�?�B�V�tJ�H���aFh�H��|?�7�zx�%A�Q��ˢ�O(|��s ����ǉ,��qm&Z##2E�&˸�v�����0H"PT�bWl�4>D��2��:���'@��,l���9��je�K,m�ی��0����Ҵ���"2���1��&I?M��ľ��w1���R����*��wZ���mj:=�e%��nr&�:�3=k����)��@��r�z8i�6?�'v��p�=�i�$�zA�r�}�ƣ�_�b+���/�ƒ��j�=(��a�i�:a$�ZȐ7����i����|ka��(7-��� FϱA	��0�#9��:pq� ˸����dv�:�f�0�td��PI7J���ph�s��d�>Kt�gn�P՝�_�I��A�C.}��*���>N�%2��M	�za`d=DG�[g��G�eD�}�z�S;Q%��0\(��"G�Z۝�yoI���B^{l�

�a�PS��
=r�#Y��ւ���/s;�u�2��Yk9�/oH��܊V)]/��Ϗ�s�$��w��jk��O��0���
����H��b��6B��L�peo����Wu'n���"�0�!��p1WI@��F�H�p��|�^�C�	n�����P�C=����=b@e�	�����̀�5���.��r��:�=!�ttq.h�������k��3��p��'D>?�ԩ{�i"3����uZ����H��!B�Of(���d(!r{����i�	^������N���X�2T׷��ā�I1ƅm�8�7���^cc}�1��L�����6�b0E|������غ�!�Cd�!"v��5l�߃������9h�1��f?�ݯ�*�o�4�ri�x��
М��J�`��վ/�RR�Q
G�V����(+p����{NF�I:�y-TW���¤t�?���H|4Di��$o	�TC\U�:m�@���e��`��A�Q�dR*F�"[���������3n����å}��G#��N�?!U��X���Of8��\�\�,�V�UҶ���0e�w�s�f���v�YC�;��\]��q��	���S���P���z|��IM{��Q3*���s��2���U�٬�1\e�<����7p8�	��d�v���Ғ��B���k��JO��W��o�ԑ>
�������J"衒�������-�p
w�^�8�E�N�����'3d-V�'|uD7s��*!g1w�9%\���OūL�$]w-X�	� ��3p��@^&�i?.Yx&�P=�ԈX���)(eT��V\[��E�O�͂��Sc���zqǣ@�s_��`QTR-
��&\���a"�Y9��N��/������6���]���]��!�҉F�y��ki�~�e�W


���8����a8����|�u�&�ے��BcuAN��T.��[�'5�z����lLk[�VoC0'S��}���ƻ1�,���n�-'���E�!��\�et%����*���۶��f 75���t-��`Ύ�_�pE�i�{{����������W)q^���4v)��fp�Iҕ	��r�9v�9����i7]�u׊4������3'����l�3[��RuQ4��	
�l��O�X��~`ŵk��������_x�sB���g�4�L����mY�.z0&����(��̀��J_-6X���Yi.������y$+�Oi�.U2�1�'b�y`;f���a��Y$��"�h����`�x�p�����>ڔJ�gr�	�V��i��u�����²�,_�ls�=�Q�Yh��g])7|���ڬ%��z*�E�' �a��gp�)=io�O�>7�g;_'��H��Y����Q��ˀT�~bo�Y���\�7I���syr!;�l����۵���va�qn�����+�*���Hk0Y@���L�ȳ&e�ԹC?���͖|�����$zRF�9Z�\�@��j�X�gR��8),gv�~��`"r���\�zu��	�w�0����%D����
��vC���M}&voH�6�Q�rUض
��*9IUҊxz!r�����t{��%�l0�ͥ���7w����4��}O�Ps��ko�m�С:�q��n`�^���d�o��i.��8蠘q1��!c�v@�7O��U)tq�:��ꐈD���Ns�w����Ѣ��k_������:�7ko�D����=�ph9?�M'�0 6��/�W_߶Ҩe��!
n�1�����~{ z���V8�'~��4c�X��y���Sw{Qҹ!��ۼ�����Y�H�����)o�Gڳ&�@y(�U�W�73Q�x2&	D����_�����4�5�H�O�!�t@����d��v񷌉y��-[��ԷK�z�I�ɮ��^���9l������`���-t�A8tD��� ��T~m����J�q\�]�&}���e\��*TUKPYR�B��+,z��3�c{��ˮ����4o�1���b&�':0�x�3�T&��8��+Drv�n�(����u,�sS�'K��"��d���(xE�R��5�JdMs�7�"��|�!�T``��oM�T�gv6`��2`����l�c@k��I��S?����� ���˨���\���I	7_!A��c���,�Qe�f���c�HTuw���*�UaO��ѧ�D��C�/7���)EA{�&U�������Ë��,��07�y��x��#������mK3�5�%��Em�v�φ9Ui��
�K�����pe���*�G�!�[1���E��6��95>Vɼ��(q$����'~�/-Y��O��;C4�&.��^��G�aL�w�i-�)/��R���^�mz�~R�e&��k��=`�PFbE�ȃ��xƦ�����{�Ho0*��V]IL|�%N�6�큸�-k������z��@��F���K*��0 ��å�4��-Fk�Wm'��H�Mh�̐�	h�_�1���ۧ�W�*�_j��|�S�â�r��2\�%כ⸌�F������"C	���r��DR��fQ�{��I|�KBɅ���^���j�|
-�Nw�K<�8���E@�W�#i&c��}H"��k��h.�Vγ���WA�XP֐���h'A�W��9+�Q��X�� b��9Kz�۟t�7��_��p�����0o��d�XlxVHYEB    fa00    1500J�\*��#��/8�~������$4H�w���ڰ#I��e�!��
o�*n���A.�Ԥ@���Ns b�ZO~�B�$�gHJ��%cCH����.�B)u���*HV���'�$٩8��j��֔�-*��C�6٣]�)!��,SfER������B(�4X$f�[���>FcD�[�ٻ�@	�Z�*[S��̔�W�{,���˘��<�`��?�-ʰ���{�NټŒ(��r�}rNy�=�3�Xc�t��nL+{��)|,���7s}tPv��Ʈ@�v|7t���LE��&!����G�#�
��F7/4t�➊� m`�J��k�ȫ�����#�4��y��;؛�!�o����t����"�b�8@(����Mv�f^g�ڬ]��+����YI��_� o���ʚV8d)΍��:kZ|3d���r�(�J�@�t��g��l�C��4WM��/�D�:ӛ#2ug�5�=��A�AK�˹�mo8\�[aD�ѿ;��d��THy��g2�ǶU�� E���c�F�BbP
����A�?��5ۦ����ݲ���>7�֡k���u:�R���^�՚Y-�7<S��j��O�_�M�T�(���z���>Iz���O�9ɩ�Z��Ҫ=%j6
�C1�S����C8�Y?!h[��Mw��ibt����S��@L?���<l�ؚ�
Ԧ��L�YX��
�Q]u@��FF��K"�o̯�ޝ�t�M�i��?��Z�ϸ�فG]y��&����z�}��W��R�>��ɈwC������ds���k�~#$���������b�5��Xm�]a�^��ϾE�s>�����Ɇ	��r/ 7"on�P�;�錓C�{,G� ���=�G�Tr����k�j3=�JO=4X����Qx���1��%i%�ݓ�.�o�jj@���R;e�^�M��N�EX�Bp�0L���Z\�8աE΄�h�ۑ�GNwI:?�=~n�Y�I����}��&����e=�z^�wf�%:��pVFs8�~sK���-6�+����d5�ӬC���'�d�R�B1�s��RH���Q�BVH���'a��X��>+eT��3�� �,<�)���-��z�X��u�n~�w������
�e�KG�ʍ�4M�z�������������q̇�5vy� ��X��c	�����$S�B=h6
��9H�BG`N�c����uS?}7;�� E�x��C~,Y!�[��O��Ͼ8mF�V�55$NW-b��,�|�c�T�D"͙��N��՗��T�]UO�w7����o��,}�{-!"����,���z�z]�O9@#��o��Eu^��q������k�0�ԁ�ae���8�/�.�̵=\h?z�-k��$3�r�5�p����x3Cit���#�����Sm)k^p����A[>����N�{baS�.�����p����`�:���Z=Hkj��xb��R�,j�f�u�o�\�� =nO����cA�0��C����*W)�#�j؜	�i���tA�0�\iVXд�9.��Q'��/R�T��2ߖ���l��(�� �cN��2Gޟ��l:^핵i���h4����Ӿ�&���o��d�b�sM���)2�׌ex�(?�^N�M1�F��4p�?~@_�Nb΋= ���j7���"�-Z��-��}�X2�G���a֕^�(֧����G�k�"O&���Kl	E�GQ������x�H�<�ha�L+�Sv���B��������l�A�挂ƚ����<�WW�#������H^@������a�`�� �J���r�����0�)p�rq�׏x19N�eb����a?��:�ک��v��[ٳ4;eS� dfzQ�����%:��tT04�������.>���cό:Y��_�����2v�U�F@�*��_�Y��������-���&�1]#�ؔ5�f�U�:��`�Ǭ���>��B���	Y䎃��V��o�+ ���5;�f�Ri���<�U@B�U*��u�h�+k���y�1�C7����������v&�Xϫ"+���s��Ț���s��t�w�4П��$���ҡ�4�A���H��aNL�H�c�L���wF�`�>7]�/�?g���7(�l�Cή�Ƴaf{��! j�/t����4�J�$ ִ	�˿0�/�#�t�|��T����%릈�xPާ�	:�:����'Kq��ېX:sh�������w��2[E>���'��VU-��c���c	��!B?ƞAt���ͫP�^�����"�y�6s���u����p9)ڗX�_,m���(&�0��g��jޝ׹e���Mj�k#�"rȽ�dN9r}��h6X�,�P7W<7`�y�Ry4}ԞO��A}�TFI���e=���*r��G!-���<�1F������Ȓj ��bq��<ք�����h����S��fq\�eu�H����I��𸔣�~F��s��ӽs�����'��L��ğ��ʆ�ڷo�����3�T9D@5�i9H۬[\uR%0"�x�f��dk����2D5{�=�k䥼l�lEef� �d�6�o����fk����~Z��&��䑷G���a=i���9��K�ȧT	��v>�bD-���.���|jw�Ƭ8�Bsnt&Ֆ�!��������^��OA�ɔ������nͤ�8�REБ�_��_g�R�E4�����&�
�H�f&H2f��I�v�m��Z��C��R7^��=ԮHPz� �F�2/�1�*���\Oh_�9��7B&��Z�+�������i������NDM�9K��l-7f��D�*R�^|�Œ~�;�zH_������8��7���r��z��	��	��o��
�+�Ѷ6�����^��$���c�<Q�(8R������z������{�63�\�~���%���SL�K	H?��Ԭb�h<e�~�Ĳ��]*�}�	�1q+^5��h���N@�J":�q?(��(��yUVرL��utC���n;��i�)���79�Mn.c��2��6P ?���u�����`�b(Ֆ��r��R޻V@�����ka�t͇q���VF�����]�nQ����P��O�p��n%{��'��(��ʾ�R��>��/�ڊ�nqa�="�2w��T&F�`.������mJ6�+J+�~�)�����~�T=���L0��l������l�G��o�ht��˔e@ҩ���3��Ut$�x.�Co��`�2ߗp4�v��
��~�ʑb�L{sQ�� �- 8�<e���E>�-a4�fmq�(�N���� ����,dLh�:���d�|�t�����N��5��.��./�9��1J�H� .�e�}4S�w����&�� �w��&;X�G��>e
 �|��!��v�P4}p�3M���i��M�zUR�� ���DV��6�bQ��ad+9k[dʂz���m�!JJ�I��ԙ����P��n}�#��G���00�����ep8���,�߀ �a�����!<AQl3eO]�0�YϤV�l�P��p�,�A��D�Z�R�Pi���3Vռ�\1� �_\��Y��*���-���0�b-d*���x�MV�|6y���/�ȀV�9γ�´�v��&��bg���*�id\�%����&���V��Ұx[���x�,�\����S�{vf���� �I�=;�.d���H��;zqv�璲���ߡ�-���P8��3Y����?���BMA8��L��,+���f&�g���Ȁ4!7�2m�X��-�J��~�ћ�jg�9��	I���$kt&O�4�@ �!"⥆�#s�����:�Bq.P
 ��a�-$�G�$�d]����Ti�:��0("�:���μ��hY���I{�d} ��(c��N��q���h3^�	w$f�X�S�t���h�U�;Y�C������a�ݢQଢ଼ʗK�)䕎Ns�X�d2�ʌ �������<ٳ����E^~���e�<��m��trwi �B�����5AUط�$Iy�BT��4F0D�/�&�j��~��\������#���$�E?0V"��5�R�^K�<�iB�N1i�����۪[+�+@�"@S ����yeҕ�i]~�����ПC��2���-�8�U�,��l3#�J�hjzf]Ԉ��W�,�u��,
,A BY㾰L��G�"�S���b�W!�`����(��c����9ʡ�J,����k�n6�ipD}-���L��/G��ב�r�S��,�Wʍ@�'gVW��`.��HE���LN+�}t�|���koV䶼�-��ot9��B6MՑ�J�3�J�59NW����6?�@�_���Ν��\�P�[D��ǰ�:����n�L��=$�	C}���;��zֆ� ���
����V����>x+��@��T����	%�5�D�\�,@X�|�yC|���ۥm�b�<����vU�o�H{[/1G�����4�I+o�e?j��/��;��t������/E�d+|�,9��BжATv�44�f��	d�_5~n�MO��G�u�B�(x�s��p��j�1fd9���z�`�M���(��^�l�M,p�"����������꼲�����&���˾��mQH��Ǣ�@P<��N��v����(`2z�$�jLϼ=�#ݤ�e�t�������^��9���� i r5z��΢ʷ�ud�'GI���RQ�	��^"%̘;L����}b�w�$k����LH�����w�IQ���_0*흂���04���KTZ�)nA��.�#㢐�E4��(��Jm$���^��%t\�����@U�43��
�@�s������/���/l\1焔v�GCA|��t��whFJ��v*)�`JvEc�4$�c[,�λ�ǂ֎�˭��Y;&��d7q|p�Co�0�N����Mg���W��rp�eJ���J���;S�)
�틀Q�����0'mK�6\�$v�i��<�����$�Ne���m��>q������ߔ��i�U�����{ �t��]h�#ɼ���� %�B˩Z�-�;w�u�竬ș�npY������`�y1[�l�t��I%��B������I�o;��i�T��%Mo2F:���x�S/�į�_]WfdW����e�\|!7�c_K�Ι�S|lz�OC[���2���ʝ'W�wKd�ښ�R�Dh_[h�:�y�i_zB�rb�]�?%<^q(1!6�$�R �1'Tk�]$롒��QV��-���<�J��^>�8�4�XlxVHYEB    fa00    16c0��(���aʖ�~��
�J	.xo��:��8D}���&[��x�w�܂X1����߯�a,�Ǝ�o*̆Y�H')HW�"qb�#.a检q�-�X<G	�Ѐ��V�ݙ=�4�d)ڤa�
Բ��ا ���f��AG�	C�A�q�����Z�G�_3Y7n�WY���]c�i��3�/�g�k�׶!WSdx��[T�b�7(�W?�#���%x�,�	��_�P`l/����LՁ��V1�c���A�%��z��l�"�m6\���C���2%1?�<]S�ʹ5�	�� Q�9�3Zd>e�=ѻb��O����3E'�,�T���~0"�{Euzq��Ў^=��3 �27�Z�X��X0.௫��[m����	���_�P_&��%�Z��Y��?�|�t�*Ϗ������f]���g� }'�F!��S��D~���Ţ6,K�eGr�+)�!��l������@��L$̌I��X�f}ܬ��cy���!�B�����6�6��m,�up�3�Ή���G���\��Y��WP��8d�x1!���ʀc�߬d�dۂ��$v���r�y��uN*K�hC� /"$�hǭ�K�7�?|@�_���xcY��?;�!U}j����CFp>m�����M�(���>/������)����t�׋��lR��H��Q�6�ҠWkC���n���]��8(���fۓH͔6�E/�K�=K�h���Dm�T�j� k�?�kq���_A�Bfz��k�@^9�)PYX�䦴F�<v,��]G��@�����2��+�ڷр-]�sH^#VcΏ���m�`� ݞP��}L��pA�Ul����4%���8�cS���2�넏a�i:8�/��u't֯�8�0{9nM1_9�cD1Z�D��豈�i�I����]���܎��Ź�t��B������c���.��z�!� �\j��g�L�ʟ�/L4�#���rV>�z�&�BX
�r��B�!2�m��t2�eQ���Ӥi�6'&*��L.���ә4}>���4ģ �A��\�s2�@׆��(�z�#5�#cDƐ�eҊq$@���>��9b
;*,{a
�V�Į������߆��uH�􉶔�Yd�?�8����&�2 5���	K�����d��\���&j��}(Z���9��f6}�Z��9lx�%4Y`(�}.��L�J	P�$��	si��x�PL�����������Nxd�m�+mn؀e�{���^��ͤ�������2�&t�~�ɇ��s�#���f��]ݵ��[bg^.���I�ށŽ)߃wZ�`@�3�$�>Q�Oɬ��	�8x�=d8�ST �����@��YHi�yrB�q��3f���� �-���L��d볻��/�w��9�p/ܟ$�DL���͐"�aX⣨����~�:F[$�u��(,�W
�Ci�2������!����J�Z[���2h@X��]�_d�uMJ�a�.]�JDq��}�����L]ꗶ}ʗ�,��5P�M�����Ap^���B	w�{9�;^
��c �Oh��;�&�3-�s����%��3.�li�)U�,Jz�G��9��[����ܑ±��&g��������.l�VΙ�Jv���95a0����:*Rjd�d���Ixq}&�Z{��X�+�9�	�bt���P�A�j�<�Up�~3�4�&���6A1u��M$׹nӒ�8���
th�ʵ�{=v�8�(;��}#�)N�K�Ϻ���zoZdD��m 73$��k
\y���Jfs�����0D ,�������zH�"/}z��R9R�k�9�^��3���pd@�����hйuG��)+�c3��iBV���.
����k%����"Ѱ�Ѷ�b�Zܩ��4JQ��:�b5��A�Fy��a�Ϭ9Q*��Dҝ��%c5�}�jߝ������1������=<�u���"�i�JcdOs�(���X�cpf��ǷOvt���1~B8���+Y�؁�I� ��6W�T��}+h�8��l�ky�e�F�.m�rB�dX���ښLF� 1�/D�ī�!�S���Й����=����
�Q�LV&��);��3����R�B�4,C�Y�[|�� ��b����v�j2y�q�����eF:��0�i7�0cԴڒ���xȩ+
�*RȜL�4S�$�[�8��.sђ�2J��ݴ�~o������(tx��U�J��:o[��>�W%���c��)&�n�1'��R#c[x���N#dr�k�{}c�!���5C�#�c�撨t�o�Y�]���{<2n�m��]�׼f>��
�����u����F�ד��%��hx�͆�m�!��U *������e���ndY]_�D�f���[���IG��,��0������x�x���D 2�5b9�'C0�t)�ౘtUR�ͽA�X{7�^���5q!�w� ��*d���X/�[�Xۼ����6Pּ�v���b�������m��-3�} }r|؉��W�C\5���B6L`�'L��rj�색�����.T��㍑�4�Ӛ�G�^j�e0��9=� �M/qw,���|;��>��J��/�:�'E�D�:Yk���a�<�lwt_��+�y�_M�(�?��e]����L�T�g3ה�ƨ�s[dit�2k�Ղ�g���Ɠ�b��-��k��1P3'��]��%�����~���7OPw��	��7&�m�.��D�9�àͭ��}�/x/���o�Ј��efn1}��\���1�:M�`�{/�"��^Usu���l��?�#*�<.��)�k�w�,�K�]))��^R҄1�Ҟ���P�N�wYgD9�)�y�&	;*���ւ����Qwrԧ����i�~O��v0Q�m.��A��.HC �x�5��^���Qd�#YN�+Pd=�3�n)�,��69O�p����6ޒo���&���-����+���7׳4^��XIO�W[b5����Q�m,#^\���x9fw��*�����&�����?��'��I4��[%9W.б3�<x�,���l�N~D#�L}��"���%��)�,�!�N���W���Q��?m�]>s�;p�!�X7s+��u�2��S���Yr�wC�n�����O��e�wF��ܰo'ۉ�	�O����e&�z��v�"�k՛�����w�(�?R���O��\b?Ǩ��,�f�3���V�N`%���3Pr��:�$Yt) ��M��4U���BC@`w9MT_�
�c�⎓g���3R	a�1�O���B,|��͠�8i�ai��N�De��C1��|@T(K����/�B��uJM*X��X�_'�yɣ�k_�r�[�~�Snw�>�|x�B�����zr�x��§��&��b.���i�������SpP\ ���O�>C>%@���Ɋ�4���m`t��)�P9%���oj�!㚫���,�fC�Z�#�9�t�V����U3���zzÂ����r!#'j��V'I��Ě�
!�ßx���}��m��Gڑn4�Ҹ��0���P`���_�k��%�b�_�l?�ˠhح��NtFf��x^��K,^ݥ��f��"~Ir9Ś���R��M1�8��|��M��YgI��Yſ����?N��vDwo��u�c�t_Wb�k��̛���Z�v�5���ҭ@�)��'r� r~Z�`�4O:$z��eT�� �og� [�F�N�689����b�5��ʜĠ�)L��sq T��|9��w��Q�٢5��i��^����-���7�t�ۼn�Z��¤ߘ���\��a*H������$^���k&�������V��$}�۟Qy�ga��b��h�\�1��,��O�yz����g�m���PR������@�'�$�eu�� �	�z��[)�M��&ѕ���ȹ���?��,�|+�!�o/6%��-�T��ۢ#ʰ`���������y�ӥ�FKɱ�-�2%�*�l1�z,)%�1�d���)V�v�~ `���X���8qWx.省gF��9�QǙdۼ4�nv��yɥ��;� q��o�wy�s�4NB>g��;�9xhCW��	�R[�Z�o��6�>4}��fxl-�&q涂������RD���N�����!`߱����,GC�W��-8�H��F�7˨OiJ����������r1��5m%a4�X%����b�K������o�e
�mg�컯�S
g�5�g��Nv�cO��Lӗ%��.�"څ�ni(�ȣy�[�Y�����Gi,U�*
u!�0�<��{hɉ��bM��3���z����E�ۯH���M'T�.SI2�?��?�?��	�[2Y>0�������l�h����NҺ�>�1�É9�\r�C�j8�0�~}�Ȧ7ɊW�F�b�H�k_��/������=�NJ%�{:�-����ެ�4靪~�)l���n+ш��x������h��x�S;�YŻ,%����-��7�ʽ'jj�u�	�T�o5v7ם�S"���!͊z��60�6��ǣy��uB��Tis\"�Fvg���DU�q~m'xX��_�|KY�G�o��"��J�T�ѽQVf���HD�B��vz�7AW{���k
�
��"ޗ)Ή��y�m-u!&*ˆl���.���F�U��.����`��&��Kned�?M�qw<����}�0����-m�Ć�e�[��W�'�}p�S��%�*rq�͘]lG�CZ�����D���-'׹�&&ϵ`S�AltG���0#}����~@��'���]�}���i]�����uB���7�)ey��78��(��_�hŚ�4%)��IRGc/���/�I�x��ը;��o^}����S�dm��C	p�����[RS�2*W�P�gY졭�b�QC�xm�������2��y���.G#��v +ѕx��0�y6ǖ��Z��v����d�;�F�:9��_���!k�����d=q�4�U�0E���:{�'W���������&*�-�m�P�r���~R�/z�F����k�ߦF���$g���iz0DuCH��6��F�!�xjy"yCG�I���X<�v��,. �H��kƃ�c��{�Z�����%�qh����Kc�pI�˲��K�{�B���Nȣ�Z��[~7s|sKѳ�{J��떃^P�R�c�p�K�)�U�`���"���Z���dW'���7�\}��[ፒp(�ȑ4���I
S,R�׾��Y���u�Ε	=�=
J&ƹ��4�e�}�_�����,�"�MX5�&��쟾�9�ڐ�g�{"�{�R��r$I"��#��S������i�8iM�g����q�Y��:�~�E����'5��(U�z����R�t��M��I#�]��mr��py�6���S��{+��`tG�����\�X��̹0I]O*#��{��J<�NĦ�����=�|kC���=E�	]֑2�!��h���a�L4h}]�����o&Z��q�)\r9O�X�M��ͭA�Ħ��mK�ӿ>��*�zcP�}�f�c'4�Ԏ��2V�S,n�=4�Q�Z�Rqz`�ŴA���i�ej�����1�(߬q���=46��^���?�1�qk�������y�`{�3H ��%������M��Zov2�o����	���b�:Pph@�o�/��RN�Z������?Y��R�Ζz��Ź�@�r�äNK�׼��׷�u��z�O��}QfB(�w ��2�t=�t��@9XlxVHYEB    fa00    1740P{&:����yL�M?����`��s�2uk�����S�����i_z��j� �8���#�[����B��f��t�%���'�#�zM��`��L�r#�)~��PLT$�$^�݌+_��/��օ��Y�L����,�:�qg�P�El��5�M�v�4���~�yHK�̴|���H@�Py旗�δ�On��ԫ��P
˔@c���o��hs��N�V���:�!o_��d�v��8Y0j�=$���獝	T�3�ɪk����(
���r~֬r0}s���9�� �1*8��L�
��c9�A#��-��S�K���Z�w��X�@���X$�;��J_����<���(vc]�Z�����@�Wq�:��5æKl��5` �S%��=�i,���&���ؠ��� ��(�x4����H L�4z���-�M	[9���+^?j"�͏�0̥��{!�M|���b��h�n���j��
F�[����ײV�{Y�c�$"r�y�rO�U춥z��̃ړ�f7Q�C���"/7�+jǤ5��A�M�X�A���\%�fǄ�c%���hu��O����$��@�l�@Q�&6j�dHbj�\��L'��e�p���#
�۽�^�d�"��u*d~x������bX��-*'
O�����Kǖ��g� z�����@��l�OG�K?��a������>&��z{�%���O��J�!MT�\m8�^�a�>)O��'[T�EG�qń�������t��&,���s�F@ѢB�XL^J
r|cĤt�qJ�(+���|�����	���-J�N��
U4��ë��)���FP��T5��'Jq�5ٯ�3�Ϥ��i���1D� vؐ�̈ǳ���8ZG���͈b���m�h�r6b9 h~9+��&f��J��)]y�T��X�_�\���k���>������R��h&>CQ�	�2�[�ca����R�B�2+e�\�O�RB+��M�$�RS�̳$�m�����s%�s�39�>�Ģ|F�z{�H3�ͳ�tn�q�Ȼ˸�!�e=�����eA@��I�Сe �C�>N�?�0$�u�A�ڊ����>\X+Sp�����ί=�8 ����r�`��Mv���Z�@Q��@��w4�y	r��׆�( �e@s��7��fXt��s�8�?w�a��Ҳ/���E=�s8�59^��R�O�^@�!�y�S���/�zj�����5��/?�E�[Ņ�;�a��0Mg��ˠ����lG�U��h�SW�����f��3�l��xg�4�q��#�[��^�� ��bio�T�Km�\4�#��e,b�(_� R����H^V�5{n�{�U�����0n�{≝<�!v�0d��z(=�~��A��=�,�j*�u�LǿLR+��2R�y�]E�X���̥aB�dZ���8u+]f����c��_��� kn�G�a%����}�^�WA���d����mi��`9���袝�<�í��F� �^tX�������a�����5<� 9��������)Ԍi䳝g`,��#�
�aN苷6ZF�V�����4�O��|���a�7�W�_E}��H���N����L#�>�AJ�+d�Ro`�~w[�BZ~�kt�~U�p)L!,�W�*�`��/���C��_�@HK�������maHjY��0 ܫzK0@��v��/5s"/$wj]���L_�<.���bfՉ�����F~2�z�Ǝ��:Ǉ�25g�r�	����`4�J���6�V������q��nB�.�6Y��v�mW^S.R��V��0V�<��ո�K;�t "�j@	�"��04H!��`���[6Ab��%�SU8En�+)��y0���J���fe�S����m���E`����C��f�n��^d1`-�p�Kh�ׯ���*P1���ȠO�� ��OH��xT%��Vܞ��a�W_��%ܸ���rX%gI����U㘎��pŏ~�<��U�&��rAW2P$0��갩	�������?H���f'ukiސ�{B�v�h���`��4����$Rr��lk���2�$�Cf`��� �(�J(X��4N-�JI vQ-E"��e��-�$v
Z/��O�C���K�Y���� �	���<���]W֕\���, �湮u!�{�qY��5_ym�(��?�g��&�>b��4b��~Uu��`;�88r��zy#��>��K�2|=5�����z��&|(��2�v0Q��zS��,1Q��+9�R=nI�F��HMO8��gbw���Fެ��4�;-��3K���P�����1�r��,��nC�h�)��fZX����''����$"I<�J�x!0�f܉�z��}�����@��}��4�Ǽ���ْ@�.5Eo&���p�l}�,t��E��PA�B�b�F$-rC�!�2&:Ȳ.��x���&"n����Q*Z>��M<S�6ր*Q�pzŅ���,"]������47,��gVZ+}?ѩ���
`�_�:.]0І/�#�q���y�\{}��t=��`��A� F�¹�=����If_p?����&j���yyS��٭�rf�:R?q(��l���y�Qנ6�d}���(e���2I��1v,`.�AI�Z�\~�vő¥?\]��i��J��V�e�Zc�A�e�>�:*����1��\�NI3Ui�r8��!��ώ.�N�Cqh�d2��6�+�}T���z��_�)� Z޶{p��j�A��H�u�s�>���}V�Ã�_��/�:��r��$+bJȆ�p.�@�=Y��%�4j�}d$��H��Cu�n+p�m�e��9�����.yh����]l�q�e���S�+#D�%O��R�foHY++�3�m�r�?���K�^���x�^�B"�`����.n(���r���PlGu�)���+�u����9�$6�^E &|�#�	)55A������+Y�|���L^�C5l����HtRAFM$D�7����6��kԐ�ڼ���O���&��8��G(�����P�+:�&w':O`s�i�E3A�_ �*4"DrpҪ�=�pF���6mȖg~��ˏ�/g�%=�]2�L�����7���<P�~U늒g_C!Y���.�]�hN�
�L1�F)����:�z8��L�C�Pi��/KC,��-�Ł�-�H�h5�	� r��Ƨ��#ή�G�'B�.�ʾے�G�K�xeX�$H;�UQ��cx���j��R�9k*�|ȏ;���e�Ek�ۙ�4cW�J0�c���#��̶Yꣴ�<�16�O�[g�y�6�grd�?�����~0��= ��8&�ہS'�mg37��}#`�(�P_���es���Qǯ?J����E����E�ᆼ���}:Ϊ;���v�:Pr�8&�Ht���Jn��+Ý�C���Ĕ��<��)agM��X\�����Hs�)P�A �@�(hLP��Y�&�;�Lȼ��f�\��ƋZ�I��]��hu%�`�!�z�@Ƌ�n�3&\���2�t��ّ<��6�^����i��,�a�͂�&�Y�[�]��{�NT�2I�f���P$hO�-}���d�E�1�&f�:6��o�����'��bg��y��߽Xk���o8�]�����9.�K2��ϴ��+Z����%���JK����{�7yu*�]���.��8K�2���^�H k-b]+˴9I&Cl�.*e8����)fat�I�������9��B�̒�Wщ��5�����iլ(-��x�djD��0��ɻ�w��b�Dץ><P��@ּD;A{�z�;�w���lL��M�)qu@��7��K
�k��r���j�7-f�_7!�(I�k�����_U^�=��(�ݵ����V�^��j6�U�3�f��7Ry1.�ZA���~����7�Z�o��h��>���\\���3������6��J���a���?�r�J�o|���®è��@�=9	��esHv��x��T�� �AG���ye$$^�ix�,[i��	ӿ�8�Ԇd�&�@�΅_�dջ#H<���Z�I*`�������=�dh�������Ar�*����A�TȠ�z��)�q��ES�\2Ιj�����a��JGy=3��aK�e��9�>M�JP��ܜ�>e�b!:t.�S�궍L�z�")��u_�>E��J�8�{"����s�;�o�	�U���U�?ʌ2��#�c�s����n7�7|����T��I���:ѷ+�o���j��3]c��$@�At��h��,l$9�D1g��*�nO�5�[tt�2��!��ͨ�xTƤ�we�E�P�s��\�N��nb+�v����6�%��8�ǔx��;�r��h�X�i��]�]/�����d{~B]������^�|�<y��ݺF��=�U�����x���'��}�Q�\Q���?Wy{W����ҁ��ꄄߚ�<]�oQ!�^��C2��K7�>�*H��Wǫz˧�Vl"%[p+�1h�_{�ͣD�E����ن����f��u��]@-ՐX~ g��`��$����՜��X�B��:i��M� eQd�(������
x��zU��x}4�� G������;��Ӊ4o��FE�A�|�IJ7���}���\W��C������w��^�c�`��X����^�:���p��.�eiHm���Ra��-|�C���&�-��bP��I����q]@Ӎ:�ѭC�ސA]�SjhB�G���>1%�X_X���F��B��4<Ѡ�&a���I.��"�Vg&� -ݠ�lC�b��,�E���ݐ�X.hG�#Z@�ԡ9���t�H2�m���������g
'D��(˹�`WP �)'|r�|H��[�S�Cq���"����Wk�
���y{cU�C�2l%2y�Zݶ2?�2��g���IT���N��V���t��!<�(�cҺ�#3�����������TE�S��=A���|��o�Hi��b6ݟ��O��Y!�)@��]($Q5��n�wb@�ðȦ޸���t��p�D� TA��(?�����������Ϸ��D������L�+�
����~4�ƫ%3)�tq}U��c�0�)(c��@��<���ۀEK�B�L����@�K�>l�*���#`Zko�6��l����ԑ�ih���������҈�'��Γ�Q�&�$����UL���J|3.S�Fb�x�G�tz*�d�0⥴�p�Z�L�R=����K����DE� ���Ω�<���'�E�[l@�~��RBt�l7��B�v%�|�V]���O�Yx����	��![�aZ��J���ǔr��PӖ�g�ɘ��%�JC=`�'��e�#[��\�U�3��2&���&�8V!e2F@� �p�`R���,0�t��d��ʯӮ�pO��C�JV�_%x<`X�G��\�J=;T��lm�G�@����e;P���\�]a^P��w��x�OIe�)�{�i\����J��|�i��Z�]�:����ZPp���kL��|
eˡR�z�Qnz+ ���]8��/�P�~�A�B������
"JӗA��߯l��Y?_	�Xn�@C�v5kퟯ-�,L�^�~Qf�G�,��|	��l��\C��oOzu���E^7��ˍ�4mP\յ!X���j}�n܍�s�íΐ@��_��(J�y����-�kf �_v��ȏC��95t�?D�!q/!���9����H��H�JÖ�$qS���/��!�_�v^A0c5��?�{��TX�aJ�Q'�>K2��B�^19�LQ�(7�j����� 3��{�d��F��f7f���ҝב���w4��
�T+���;����Y{��G��XlxVHYEB    bf14     c60��l���n�R�����c��n#�J�ߏ�(H�\�Nоg2�!� �V�Ĕ�&�.���7
Ҏ��j�kdJޟ��UT�^�8�on�%�aD���ͳlԁo�u!Hks�;�:A S��*Fv�Xp=:�^z�"z2�g�U�!�)X�32s��զ��`_�	p�9@�P�[RG��YJ�<�<���89�P˟.����Xi&k�3u`/��΍���ڤ/8�,��\R<�}w-����߱���M�ꝼW�WC��g��E=�`.G�g!��uј��3p��y��VEDi~6���ތx��b��dյ ��T��qf�s�M�*�9�q��R���,���'�4��Y2i�R�:m�#	���n�I���JqlvD��F� ��I��X�|r�w�#�,�lN�\�s�	��X�8�M�Zf�Ү��>��.HWGQ�{�`�ƞ��m���j���*.���<D�n]�
�+]�9��=^�t�)�4 ɂ�q��Y�)���~;�#u�M	�;��n�,'������M�e���+�r�m�ם��o��<����LWeG� ��О�� �+�	�]k�/�)���\'	�*Ұ���#��U=�#�|<��tڪq@�E-E|��e;%�z�SG(Y4?V���0`%���9
V�ư
�(,q�
�-w{�����+�05���9�#�M��3��c�t+FT4���ޝ|��C]l|]���.�J1��dd�w�g�x�?Kv���PX�@Ȃ�Y�ũ�������
O�/��j�C�#������$yx0��;Py��!�����s��b�6�qk�m�!,;�s�<��w)IBǱl)[�]�9|�/yD# gp�c�T��;m\����,���I#�E�&Ԏ�<��Qt0i�3Ⱥ���Ɋ�`������S�P?:� �Ù87�cG������+L���K���M-}���e�<!�Q�*�������������rm z���r�Ԏ1���@&��F��4S'�a�ٚg�qzy�[^�
߃��"������?�0�"���64��{D�%�~(M܏6��ǿ�%�f�ٗ�E��o��r�*��w. `��FV�1��{0&B������>���ӑ���O�e��
�����A
闯M�ѨKo��H�efw�eE��eZ�n�93�o���7Q��C��iG��2E.���{�q�]˫�Y�������3(G54�����(Z2�K~)nҺV��f�#�F����H��pe����8�r9_<%�A���2X)��{�M�Es��Z�4�2~��޽�$8�x{<��׼4�@���
�����QsMI?���/hmP�7{�m.m�iLCL�8��ywf�M�@6�N�5���PeBJx� �c�m��:���>��v��˧��90X���0~uq0��lb��\��~� ����j���}����mWÍ��]o��.NW~���ɢH�����_zP[��F�!�o���Q��B��LM���#�0�Y��xm�h�������s2�J�BZ��I�s3�����Ta�k��E�m ���+[�����h״�L�3t �+�G�&����݃��8�w�$.M�������]$;u�"��U���ΩF���Zy7۝R����ȁ���~Z=Ƌ礛~e�+�~럻Uk�xG���\�Q�Wu���W�#�82pw��4�#7�ڊ��kz�rS�II�7��Rv�����������ď���|3����'ɽ�A�[/�����	.����<�in�ٜ5w�:JK�� )q���ߋ�8t���j^E����R`�g�ɝz��k��c4*�g����0)�tn�Kp8�(�$aď{��Óۄt���[�����e���>R;�K��2^���.��k�O�gz@���6��o�~5�ѕh�و&�0"t#�dR>B\��v�(���1r�!(�ǩ g`1(S��*2�?a��k\��2�!r��Y��6`Q�~�2A���/��JcM�|L�黹"����9I5`��?H��vi�KF�T�S�r	O�S�2�o+���9Y<� zD]�<̺@>û��&�gW�L0 �i����n%��y�z��ٜ����992��g��u���d,<bݳd�?�ϧ�:j*�U��	��}�=hR-ӑY�dV85f�'��I��7/�G�w��7f���Q�o9��UP����;6�F0ɗ�D��Ɛudʎܔ�e}{±4ytA�J��s����/�|r%[�L�9\�. mrᱹz�*����2���NO�!Z\�s��[����с��7�~�^nX.�u����X%"k�>�_�j(1,>z>���Y���}�[�0׉�J="d,v>@\͙�+�/��T��Gp���]N�ø4�,Rf�\E��&= ���j�����p恘�:~�	I�*�5 �$�mq�<�U����ά�Z���XQ�P�=�#��	I�������	�A>\?
�x�bwwN�}>�l��=JH�P�΍P�+��CF'�|�lTSr�2o��ڌ�����/����3�C�is"b��UpB]p�X��X?�����HS�u���ήN��?���ڞ���<1��~୮�Z��g7t��1�E��?mzR@^o&����[��{8��@��3W�KŹxn��>�^�͗��k��{Ixa�����m>��9ٹs�,��%�˞#Qk8_]���t��I=�E�Z6�%+ʱ�*��&ƕz1(��T�i�������8����"{���eE���hX&��ia �����U��xd�\��%B�)�NL����o*����<4}�)ſ�r3��־�����O@�}������%���J�4�˼��'��7��<V}J(˙����aS˓!���}��H�.[ҥ� �r��#R<�~� ����\���	=��S��0%�_G��m���a�7���"������E�s�Bk�$9��t%ť;�9dФ�����	VBS
���Oʇ�d���i��D�[o����>��P4��D����gc�l�0"�m��yj$l�o�eC��^pZ�0�zb��Ug���
kLJ���G�	$�D6g t"!Q������b�"X�x��"tՒ�D�KXR�{�;D-�"��g