XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e켅��w��Zz|L-n���ɤ�D���TD���s=X("�d2����碯���j�3��3i�J��㽺��P���������2<O�����;���s9y�@i4J��,�:�����0�upk[��u�JK��l�ʲ���I;�N]��3+��D�4?�j���]�����#{�)gYU7�!7���r~�|�0��u���5�+��J:u�ap�`�e$OF�W�=��O��1)��SR[§Đ$?��<V�@Ӑ�\Kv�5�z��9��7e��I> �����Q���?���Q*)��P�k�&���cE����<��M����z����x]�7����(�0�bs�ߙ��Si3;H����u�q�l*��/��W��ofwfL?�V����/���M��ay�)q Qq�ķ�z���z|1�a������Y!}�.���=�Fz�N3�SD�Ý��g�HV���|�VP���W�E]�TjO�?��0��|J�5SǴ���`@@oŷ������(�ӡ���(�|��mS]�c	$pA�k
lgMo�r�.��^��=95��ع���(�=�6��^�	n�/��(���	
��;}wF��C�thr��5��������W����R]@��~�]��튰NІ{~�v�]ơ����Sn6-G���pT��@(<����k�� x�A㋒�g[7*O�N����W�8�{�|FA���NNpiΦЖM�c�h��y3�#�XlxVHYEB    56d2    12a0`�}+��d����4ja����Ť^Qp�0�uy�f�Q�UY���1�����	7���w�����1i��v��6�Kg�� ��w�a'u�c�e
��n�8����puV}u�H+Z�+�|���
�!�ea	���1�Ţw6]��ᆂ"G(�Lc�0�m_S��
`���N�(	��+���~�v-&rp��N�a.�����e���
��:��)$Y��D����%Q���M��ʩF�%�3����0 �l�l����Q@��V���Y�f��V��CH$ĺ�;-��׃۝R>r�"��o�KHO|�l�3�du���g{�?m��*�M:�ƀy��C���<$T�g��l�fq��Ui��*0���Ç��>0��[����z*����L ���l&��V��PE�=!'O��0�l܌�ș#w�BtY�Q�|�d��3�v�o���m���\Q�����X����$z�w���_Ek�a^�����9_����l��.�J��j��t��f7�A�b~B�m�Rn܈��͉p�/� ��������)��������@fowZP�/��V��N��O�G���F��8�G��˰��Z�c�Y;'���y�{0d0JX�@,�+&yJx��b1�u9ӹOP�ΑN�x���>�A�$���˖�I4��i���&�����_��o
�S?K�OK_�↨O�))����<��;����zQx�.�n\�C] bH+\B����5C/�֝�4TP�zS�P��f��a��Y:��W�zC�h�ze���X<OZ��r4}�@��?���$��|X��i��i�{/����PP�	JB�a�o�\քS����L��m�����%H$ٞ6��s���+T��j��+Kj�-hϲ(�8Ul�c# o,)b���b�nb&�HJ�S3�<�9���W������	�&�kY�Jz?@8t�_|$�����ە&/_�,��Z��|���D����h+-7~��"�T�w�I��q�fnl�"{y�#_�`�	��C��_d��.��;q��-�N��k&v0A��`�#A�E:fm��>b�����ؖ�"��n���TTb��A����w]�~�Eo��E�����h��MO��",sq�W�BO\�n��7�>,^ #Ȧ��/�h�K�2p7]��I���|pY�)B��[["P���)}2�Wc�0�_�[���V��^���ܕ�����H	Jq �м8}�����"��ub+[�"E��O�֐����@�2�-��� ��0�/BƐ���:q�����QCD�fy����G�p��񃼺k�م���BU���bߩ��X���%��㟖�.�|ʫ����Ԅl #۾�����@͑�j�C�>�����gY�{"��y�{>�����^%�܀���~�Y�?4��gg���P��C:��"Ġ�2�9�|[�5�����4r�����N�}�%g01Yd�܌�ݗM��&v5
�x�zkY1����81,~sBj�U��UA���>V:�Z����'X"�w���`�q��:W�9����;F�X݈�?����d�N��C��ݗs�5��jh'A5d$��!؃]±")D5 .)�k_I9�t'wJ�H2�R�s�(4MPT��FH�0kw�*;���c�-�v(��OK�T��k����#ey�w���*ۂY����<U"��]F�ŮGȪ�ط=8Ro^���3Z���ዌ�tZ��'s��b<DP	���E��2�P�Eb���%�r�՚1�F���Fs�6y�y�^kac~w�V����;**�0[���.�bz�ÑQ��F���<�W�O�pcd��zu�HB�lvdXƸ��h��� �N�>�q^S�@�N �ү*i:$��{=���=����������w�� E��m�[d�F�2�޿��3�τ|4@�8+l�7H�e���MU�3�ƌ��z��G��xPl�~	�0F7%���(�R��d�"3�`X�H�di\7�sM�`l7�j�>8+�o���
����	�~c v�z����\�	r��x�Q'
JkwlBA�Y���'b���SqIL����Ί�A2ar���X�0�Z�6Y9��\��G��~�ԫ!"�iF�J ��bYDe��<�����XS�}0A�M	ґ����n�]���]�X��,ݼ%h2$s��\c��\�ݓ�;��@?p%��Y��_�@8�#�g2�YA+"f�9
 ��*�!#�6�ݪ|�B+�6�hݡǸi!
O����[��UA�/���z�U�	-J8C�?O��ğ|���Iim5��3g�J��LϮS+�
�I~�y�6'@�Br����`���:��gW�(�,�A�;ȥ���eYʻE�E���2Xx��%���?L2w~Y����(½��b�"@��=
(S�������2�T��FQ�X�U��(G@j���mM|�pZj��vGs��Ƙ��}�+XTt�73FPC���ܡk�"\ㅯ)�C���N���X!�N���D&��)Ӳs�����c��H�罔?y�o[������Z�>%e��:��+@�ri��x���x�p5nPGjĿ;�3{��a�hQ,և���h0�J2���!	B��k6��F����{��=uE��ӕ�:Z=ߝ� �Q��:N��B�yR���\�e�J]}��΁���4�Qnt#�o
>k�G�j9�����Ň�U�b�H�A3}���=��v�/��Hl�O	]�i�)�ۑ؇�6t��� /�0�Xγɋ���c������L15��;�l,���rg��a�����[���DB�����%�޳O��]Q�δ/2��O�����1��e�Z9�Ƌ��k��2�$����
E��/��A�z�>X����0�Jc>��|��g{OA7�G"�qu ���5b��-�p�R%މ3���w��`�{����6��a�|S��-�
k���K�������/H@P��Wx���O/Sf�o ��4
�`u�����)��ɶB졡�U��30z[���tg� �?Ի���+��T�-����K����XP 
�G�����`X7���qCD�mcâK�p�Q؁���"%ƽ�qDV˹�Ǵb����9�y����^YZ�LO2Bs,���t�����ջ<(���>cx�B(�^y�x�8��T,� Sx���X>�l^����s��l �	Rza��S�UV�33{�v���f��}w�[~ٱn��3�Tp�q�оH�>NZv^"��,�	b��4[��n��y.�"���Ox���#$��	pk	��9�Q,:�b�G��F.Q>{�3�A��N�,~����q�|��'�*$ �Gg�0mOˌ�#���%�!F�R�Rv�W�5�ɨ�y	�	6���،�`��P����b�b�R���\�����2X<p��P���C������N�lm����##��Y�C>Ž�>�dz��+�B����=��(���e(�E&���� UӸ�y��s_���v��\��܏�a�\n�3���u�Ï�8eX��QJ����fUDA��Y�bMh_����Q�i4H@�=�n���Nu�/�硵"�ڿ5���͇��Gv^�0g���-w-C�Q�Z�0�X�t�vŋ��r*��e.�?�_����H	�A�t��=l��OjCV�=�hL�_K˱kJpN�$����ȅ�π>�F�)Q���?��_򙝉B�G�V�Շ͆�k֨�#�eJ$&����������Dmߒ��V;�Ŀ��$�U��ߍp��(�Dۼb�O��r2&�i��-w�>�9~w'Z��%W����*��ܝ:��2�܌�1���Z-ZTh�����K�踔|Aڼ�ϯ~ڛ6�@�]\p۝2�FM�KT�k̚F�����&܇�Ŕ4S�>�4��z���FA��a���$L[�I���H�aڧ�};0;7��e�VП	���������J7
˜�����;<"&��Ld�n�N=�/s�3ã�6�
;��W��r�k�ő�Yn�"q(���lyuHo�9k^q-+�����N-�D����g�������y�~�HԂ# ��K��z�)M����#�V��RMC��S�%ԅ��!"����P�ÌE��h��� �ґ�K���YÄ�$��t���A�uL${��B�/N+E�[%�Ia��c5Vi�EvJZ����P�6b�J�I���T�����c�l���NW��B���]e��sU�јp���"0iB�2t��JINɣ���Ixih��Tw�|͘0��Wb<M��s����_�?��~$����l����$�7했/��[!z�X�R	}�.���V��=���d>��x�f\*<s_��B�Wg��9�_�{1�S,��n�y)O|�P�V��ת8ϔ���B~L�v��1��1c(��z\aF`�c+%0���O����:H_�ؓ)P[�Rg�r�7>Yed�4���K�f+�i��u��,��7�FJ�T���V���\��R�{�����Z����l14^xK@Z��cC��^����#LQ(�����,˚�������)����~g�i�<����O�D�M��g(JǓ��G���j)�d�Y��B����~��CQ��uo�HZ�AU��3[Ȫ�s}L�Q�[�,�A��?'�;�3�P�~`Gչ� �%>O�ԟ�i����yu "m�G�����@�6#�ەp�̭�rМ��xC4�v���#����a3��b�%�t�[/�+@M�*`t��/%q{Mm�x�8��