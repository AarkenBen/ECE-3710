XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�T��=����=$�Eș�����-��S�FS��{����~�K�I��o�2`��-+���m_���mP�$�
DT�'��~�Wv�\��D�m� 5���<�&\��S1_aGS[�S4;�>�j?�������Z��R��2<ڠ�����L����c�0�O�H[d����^�9�ǐ]}O�t�G:��`��0}�`�#H�f�Y�E[Xy�f�%���̅u��!�/Ӭ#꿄�Dڙ�n�au�?H�"\
L�g2c�!=J��q����_{�»�@'X/OdLj��~�Y��  u�;���?���Ѳ��D �$�ר6L��/�Ƞ�`��5>H���>c�ŏ��Hy��Dk��P���^~|S6g�pD�M\әAƐ� �QDzp���G^J���6-[1k��^3ٞ�Qw鋜`u�^a8 U��H���SO~Mm��rh�~TQN���N�O6o���*�Q�����{�3nF��@7�~EK X]�Z���dK�?���# ����g��7��֡����yd�׭���%'�l��d�#$/�+a�`�]�Ԋj�4�>�]����WG[�=�z{v�aV��:�ϑ�β�2�n���8y'T���������k�չH(�D�*�߈�S���K�.^�Gg���C��$�r�WڣH$���i*7qaD�7l�ko�@}#���E�5�Z,w,�x���J�Ӄ�8ZO1��HY�S��H�!�~ba����Ło�����o�'��Do���|����-q�XlxVHYEB    ea93    1880؊��eN S��ӣi�g��	�`�A(Ou|���5
f������N| �c��	��*;����+�*j@k�e��NS�*:0{������T��kC#�~y�u|N��G�_-�}n'��3CK,$��/uӗ��5�p�>t
��~�j��A���zs0衄z��c���/��vU�KN�P���덌$Bb�8�둤Ѐ���$g����h��oY�G���*[P�W�C���̃������{u�(�0z_\�,�2��[Z35O��C�^F���{��Yi䎖�8���N���𡢬l�g/�#��B�+�1��K���+�c�_I�06�%7�7В�ȵKՍ��.�1h���f��/DF�ޒ��a0�gp��t<�f�[?H���8O�f<E��j�,}\�\Q ��I��� t�,�FtP �X� ��h��#8�Op0�޿�t	��<Ƿ��o�%۫{�B�s���^݊ ��+@��5$���\C���}�����>��;bD(�������sK3����Q��Cj�ب`�l�k��8��}�8�m`�>�R��ӚZ��u�r��}ƹA�[9����HW�<�txh9en���G�~�d.�ԑ���2?4���L2������!��˪5ǽ���:�b�:���`�����`QaQ���B�\���ոS@4L��&��������N�]vt?\��C#e��~���d�١ҰO7���������o!=O�O+W�׹.X�@�y���~T�L�#b�M�*��@�
˪���l�Y>�e�q��6�-���L����`����aK�ݐG2{4��=&<���k�t�y~3��@A��<�\	ap��Hcݨ��
Y]����]R�v\<h���5\o=_/�@}+�i�H\ 	�=Q̮<�׀��q/"��UN`�v�=X�b�&��,?�th��2b����5���6y�0��0jY\%��]��=�茸�ls(l�����!IΗ��	>��p^8�I�F�����"g�\�^������l%`�^���>�eAM���7��Ve���1�C���X�Y�
���+Z�G\�D�v$���봨lq9j^A(K�I�oC��5ut�5�ʔ�=3?���+3���n��).��K���$&OK��SmJ6j�/�; G7D����tΝoH�w�|�m}�y��g�G�t1Eh8��@X9ε2�i�]��WU}��ŕh.���L��|��u7��A���c+���b"�=�Z3�vԏk��
bһ�s'�o����;��n�@a���.;�/�?�Ѣ��@��b�ɤ��¡,ʎR�p�n36���o����#1��\i���4�8������K�*�xB�:��md�uW4�{BF,�X�� ᐴ�����|�9.�����YJ�3�������I����8h�XK��U������}��#4���d�v������;���Uu������R��\��U�oQ��Y�����G�{�G�Hs��"r�b6��j��eb�DZb���
F���Um�;OWPѭ\[����BG�5�� ;�i`���TQ���肇�t�h�����l=�3��|mE�`�@��4�!�X���<�7�H'@�'�J��4�p�YA2h��D�4�����N�jpݾ�d�ӊ�����vE݋~�.<1�).P�O߬�4�
��Gp�)��BSm�K�S C(۟��7��i��6�v�S�Ms���5(�XQz4��T-^��W-������GK�a�Iy�4�2����z=7&�U�Ȏ���Èpun	:�����e�����`��1Zls5��>��kB�[���[����ta~��� ��F�Q8�2</���l�H6�3T��U���mW1��ޙ�_�����mq�۽J'h�"n���S���g��جo 2���p����f����.�� �~'���|q�Ȭ��k<��6����.�cB5w�ZCXBs�')��[U|�7���N��&K����Fϥ}�rr�pm���HW��	J}�f��^�ęg�E%���a6NɅ�T�?|#��U�'�V1<%���1�O��'��!Mn�l�voDo����RU��;�9w!S�~�YV��_=�����r7`N����%�=Ϯ/0�޶S�9��fG2�ikH6�eJyc�/,��G�����Yo!'Z�m'ƙ�6:h�#C�Գ�3��c��!^��-�BC��N���O��t(�R�N�%�O`�P����?k�4;j�R>�K�_n���� M��qI�(�7�tQ��*`�֖0�=भ�����o~P��V�/�֙�*���=���T~���d�XyP��H�Gl����n�'��-��<��"�g{>QW����W�OXd��0�{�f�5�W���J�8<{�-��_��~�pu�h���S�ZA�r� <J�~`�Y!a�	A���^�0,\D��@��R��'y� p�S9~d?z�°cŉAk���+v�'F�S�@��ӧ�=78���R���Kc.'��Z��H6�C���0ks=�W<�uQS�>tU/zF����4s��u��G��J�5������-5vʣe,�m���S^H�,���ѱp_3΅d�����ث���h��Iz�	��O[�O��q�
�|��"13�=�1�t�Z$���VOyp������a/���F����TFÛsh�/,���'o;
�?�N!��#J��_����&�A���莴��}�иC��sA�y�Ω�\��	x�Y~�Wl-�2�~���-��Ί��I�W*�P�h���u6��ZGuX����^��r'�h�ɍm�&���ua�M�U*���%:��!RM��iW�\�3`������1s�I�lZ@|[��h��Y�T���/�$S��s���h�W3_u"��DT���Q�T��S���j���}1stEŎ��fP�������Q�E]0-��;\�	$�m�wwW��( (�]� {��31��QD�k��չ��H�ZJ�V���j���T����W����L 幑�L�?.]3�bU��y�!Ǵ`8��\o@�X-��jP�=��-��h�^�V��,0aĀ�U�:�C���&���P�_��M^Ĺyl��f^6�e&�k���_:�O�ɑ���R|�v1e<���ui*�C�**r6GQ���m��k�S�} C�T����o��Nh�^����)BL�v��/I$|*FHC4�j��ʰ�)���9&1j/pR�QԸ����X��z�҇y+�D��F//�SG,���˯H{��� ,�`�
��U1�� �nE1����
"�'�V=Pf5�rԿ�S��Q�~[��ю�ݛ�Б��m�����4��v	^�&�m	q��Bπ%��W.m�>�g���!���E��.��@��\}��Q��+B���Y���U��0�-W̎4j�݈0�3��X֐���ۮ��<��7����%�4��
�G��Ѥ7DG�p�p&h@��Aҷ�11��sy%��,����wG� l���[h����<�h._����|ߜ�9f�eѺ����u� ��ܻ̼�y�F�`�S��B�W.�7@k)�ys4���>l�YL8�ǊhZ�x���/2���搫'�	�(��?���SgO���������wi ��fAץ.{Li�n��U
�_9�F�v-+��ۡJDӢ��%����V��0_!�n�R6�P@�e(���A�q�r ���p�@���ywB����j�:�_'Q��E�jJ�j!����[?�9Y	{�'�|o�ryi�B��F�S�$ϣVܒ�n��9�h��[��\�=�k��҅�tKw�q+��z� ~@���s.fv�ѵ��3ӎ�`��4�Mu�tܟ�,��7T����2�1 y	l�k�}/,�c�g2PWjr�
��K�!����L,���HiCɺ�-�:8+��:���IB��=�y���+�	�ڨ'F
vK���m���[Gw֩P�br>�lIg��nȓɅ����IM)��1������v�����b�c������%����|"y�)L`rq Y����y��7��!NܔT֓����@GOZ26��D0����5�4up��Q�"c�6G�G9DT�w���CTwF�|�xF兵�57�[�m��k���}v�-�����SV$<6{�����r}A�}���>Y���OÜ���J�d�b��e��j�z'�R����AC����/ӎ·����;2	���Y���7���H�{�i�M�>��� 2���w��{ {���2!X�E��c�|�ڹ�UW��J��1�ǯ���`ʹ�о��PUц�>�j����)��S{^�[w@�QK#�
2=[O��+���d�5����݋r5x�(�>{�9��o���(��1���g����s.فſ%�� �>�G0�X�n���tM۫�2b����aY�n�c�s��9m������xa���� %�ʿ�˫�)�O)�'�c����g�3��s/��{�kY7������Y�K��3���fj���rTCX��	"�{݊\[�
]��3^��X��ء´�>h�ʫ�SC{���
�<�y�����d0a�A�`I ;6� ��_��ۀW�y�=�l�����{��z"����Q~U4D�i�A��NI���&�w�m�b�x��߈��io�*���(�K�#zyq�ޑ/��qrUi��1%�E����+}���)uRY��b�s�_�0�H������v�Z����z�W0��pt��-b��u���n*0�H�<[��R���ނ>�>}��͵m���������u!=ɫО�<�s�+���Q~�}T�I8ѷ�V�o�j�lmz���eh��Lt!�u���9zeb�oK��75����X=�q'���Ԗu��D2��^A�� ��X��#��&m���{�qL>`�6l��l,y�(6���h�5JF���>є�La�z�&oM�1��b���!f1���]�P$_9 �$�o"���v��)�q�B���-��NuLak��2ö!�:��1"`�Ym톉���%<F�a͙kٶ��l�͉�y��s�Q��!��ѐ�|��I٢5~f�U)m���w.t�����iu7�3}'��&�>'��h�3�N�R����q�ǳ��ҡ�p�t�p"�{#�rI"
zQ�aƐ�s%�&2q6����Ρ��汞r�W1Q@�C铝3_{XzZ��xQ�H�+��'O�.�y?~��t�����ў̧��j^�!�Պ�j�NP+<��.�CuG�^8��e���a�-p�+H�y�ϓ(bN��ƸҴf4u��d��妉��O��rH֨o]�!7Jy�!��}�\���G����q�u���P�J�%1s��y��+a�G�P�����S�� �N/�"ff���=U#M���
��3�ol�G����.Y~�_�]mhʬܟ��E?s�ӆ��C\M�3}+PS��XBb 4a�6"s�iA�d,��h��E�+]�X�I��n�MgX���1��#�ͩ��w�R�a�X�W8Ӹ�[��(,A�ώ�,��@����.	�?@@`FA�űM3����e��
/�?����!�8u �f�k��|C�6N�C�[B6�H%�:�NU���B.z��g��2�N]%!0�0�\i��Ψ
��3tXOK)_R�Q04O���dP��7���_�#���
�&J��N�>�Tգ��q�_2l��n��ɹ��_\�I�o��^�"�E<ŗJ�ZJH�,)=��t?Pz��g�r󨽱.6�ϧ�л�#�^`��y��sUɊ%��C*��C<�=�g'vz]���u!�QO�Ĳ��0��-lp��˷��X��O�u(��&� �[X�Wȱiᢠ�AOY2�7��a}Oa֛i�w��5�M�[�a�~A
�f���Ji�77�2�]rHl��mIvx�����hEu�{t�%zx�)ϐ!��"���u$ho�TAq����V�t8=�o����;^c��$WL�_���^���GH�z�EL'i��i(���=⑲+'DVn�Z�y��|���m�W�sâ�° ���­��&R̮��sK��#������j3P��q32��e�u���M��g5���)���E�0��0�0����ŤEO���ݗv���i�m2xR��5bK_�c�z�Џ}��t��Jܰ�|�B�Dk���3��"I@��#�����