XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_wI�Á��	)�7�N˪����~*I���-!D����v���R���̒TWr��mrlŔt.;"F�����(��Of����75%����BN%�9p��M��:�wB֡�5�
��zFy�q���dH�!�Rĥ{��Qy���[H�Y���md�Q�J7S�N���"Ot>�k�P�AT~���[�\�ur�ԏ��8�����Ǧz���-�:c��o}��"� �u]��Cb�Gz6�b��B!Bݨ$��:�r^TLGp?�F�[b���Ԥ����e���܏g�WI�[�pMV"���p4r��?]�{��kQ��FW�&oͨo�M�儞~�Z���?��Ǝ[�55�2�D�Џ�;�]��!9[�;��y.]	A-2���A��n�M?9� �*$�r��3�Ot5+���_Æ0�W��D�Bo(���<%U���������M������@\��j$�Wb�;
�^ʫ�`���P��D?��h�o�����6�}�w�SBLA�~k4YW�3��ڣUcCD������r�
����^4�����i5+��{����-Ғ�s��=��`��+�\���'���{&��v�?]>�����3�]��ni:KY2�Qٸ��n��h���n�0>�`�s�����v^{e D�i-t4,�^	�oP��!7��肕�#I5�!+�q �C1�������Ug�H��x6f�ڊ��.���wȌ1}(=/�U�Y,F�j+ݧ�)#t	Hť�$���2�XlxVHYEB    c3e8    1d20=I����=h1}r|�9���z��^FՃDf�����!����o�c���{ʞb�'Pd>q�&#�gw�Ҍml�:]����W������'�3��ao�8	ڞ���	����x?��h�i9?l�����"R�נ���CvqnETT����׸i�p�(�+��ay�ɑ�Z?�'Ϣ ��j�(�)�ݢ?��DR��.����;�����,kG�^�a�B����������d>&����Or�<*`?����l0�k���ƨ�R���Z�;����l���Ӏ����8?_����4�Lg�\�-���)�4���=����߭$Y�зM�?!|]/�_[t�ř �f���C
�r���Š}����VQF�جi�Q]��m�d*>#��V��W�8Rt�s��Vg0M�w��/ƣ����,d����G�'�oQ���4��yr6F��$&|�\��6�_�����-\8}�J���S��%�j������)�TWh#��80��v�x�J+�#>��una�ʵ[ ��m*���҃^�C�!�x��bu���XZί���rL�I������J4�$c[��V�4^���rk����9ٱJ#���FlQ�	�j�lE�¹v�>��<��7v㛙�W@[w��9��A2�Ϟ'�����1����O�Ƴ�V�*}:��u�����p����u�i��/{Ă�Gs-?���Z8ķ㱈~ި.={d/}��U����L�\���qԣP��Yq�N��@�4����$҃�%�?�k�Jvl8�l�J�.�������{7�,_�mY�Ư�H��f2mݍ�qyJ��;�O�+�A���"J`���a��ֆ(4c��om��&�.�(�I�̊ p#�S��t��Q8�a�H��S��Ynf�(g@
�đ�jMPV
�j��EH��)�5� �����.��5	Ur����c(���~B�p�p��Q�a����t0"	���o>O�6~!a�T0Z���K�R����KjN�t��.�H����;
�o��me
T�<!�k����v�i��V)����B#H������S�2E���O�<�!�(�l�bnѲ%J[�Ny\�*H>�t`��{Uk���Ҧ8Px�^�t����%�����q�Z�Sx��)a��G(}T��G����s	J)hE\�m���tZ5C������(�)*l.h¥��跁j��
����=y�~Ў��N�g3Ò�[N/q/#��!����_
�NQ�H-�\�ڦ���XE���� ��.f5��O␆��eB���X���ˁZY�b�Ae������c"\L9��"s讫B^[��b��|I��1�����z*y�H���M�DG��jHl��i`H�U�X}����<���p<�w:*_�y&���'�`A!T�� �����e�/c9�8V5B����:�$D�>�+u}��r0�����r����S�q�ЧJw�7�m��,E7�Ӫ�a�c!i�I�)A�Zi�� ��kG�I6��Yy�A?q��ȡ��FFP҉��(���G����(�l�>��[��w��1!�{9�t�δR���Nٹj�(�����S+�tO/�H�{������V���j�A��y��@ϗ�1���t��oZN�t`�������e`�ֿ��2h����P�<1�U��G�3�v16B��љy�S���b�z_�{Κ�v�xw�"(����`I8�[��1!j��h?����E��y?&�T��~���ӹ�8��9|@�n+�p -���yM.!�+nX��*D�)��r�� �D�} \fBؾ���� bJ�F�>�ƚ�!����M}��Q&���������=�D�����]��F����@�xl���m�GV��̙u�"����(G dM����Co�a���<]6�"���G46�|@�>oQm��O��`LI��V�{��6	�;>"'�j���,{%{�h��P.�����(���~�r<�LX�����~�V1��;��N:��s~��$�o?:@������|Da��cv�i��|rc�x�n���G��T�%����a���z��Y��@|�b�j-ƽ'�a�./�����;��D�g�)h��7�*��0��T �p����M�k6�S����k� ���!O� ��
�{P�"������݊S$E-{0L^�6�ܯ�x��A#KA�z�J�c�MW/�Ŏ�8���ס���}ሮ�'��5"�`��nE@�%�R_��� o�����4�Z�dj������R���q?�,�(g�bvJ�4̀�����-���i�x�xę�3؛T��'�ϔrG@���p�V�Fy^��!��u���$����^� Z"�.�ɐ��@M��<3.�{gGn^�ͧ?��9i��%b&����w�m*�o�z�Ϩ�
��AnX�~<]|�����\oU'h�&�1�i����Ȇ6 vZ���s=�5a;qa�%������A7��a��,�-Wm��*��h��I��[~p�C����\Ot� �v�}�`�FS..URx�gN�#�FIJ�(C�o���*�K��\U7�������ϼ��q)Q�b_��4?Ъab�B+> «��Ĕb蘁p쳞S�dZ]	h��w�!�Ū�_���O«��x%>
�77�l�V������Rƙ�#.s�#�"��K���P��t�I��g���O\rl]7�M@"��|�����=D�.º�iAɆr��: g��{�ZGx~{y��i����:D+]gxH�$�2	�F�l26L��K�-����$'B�E�Dw��s�����Jˮ�GV�Z�+��i���t?Q0�8�T���l�~����@1�~G���{�k��-��~}v�W���&%���"N!��^۷R�3oZr��`}.��9��z]b�����i6�S 	PKXJ���,W#�r��_��Ny{�~{�V7��{�K�{Lb���-8���B���g�*����ؕ"�7�A>Jb��O
�}��`�*�^���n1��`^���GC.������"��B�������E�2[$_����tHA��ag3H�NT�P��s[��-�9�ם�ºH_����E}
�JS���8����NJ�E���i�[S���S�h�]!|xX��L��ݖ���К����b�$s���4:���^0���-t֑w`�����7�;@�~b�� �<i��0�&|{H���WƓE�>��0����)	.��w{?��������ˣQ6��cN �ѿ�H��N5]��T�]!X꧐/Sqr�zC��?>FC��򲷱�C���L���f��G��2<Ѫ���fk�Iφ"���0�:������&U����4i1�ʙbu�V��ߧS�lY�%���yeA�T�p[U������(���,�6�؟�9 �8��Ze�EM��<L-�'.�Ix^�߬�۝�SD�����p��4s�q�A�X1r������i�v)�%�����@�]q��{�G��籨��&�)��b��6ԉ��M�'�(������<w��7%5�Fx<�k-��BS܀��E,�����R��dh���W��*�B��cl��lǾ֗��{�*q_ �ʅް������ZⰁ�@g���%}��e�U�xT'�����x_�%�[Ιl�=�)J� ��:��Q� A����� ���M3йĤ(�of��ν�]&�'�i�"[�a��~�_�$��Ba1`�s�wٮ#����ė$�����|e9.����X�}ju��Sʳ�B�C6Є$�ʚH�)���!�N{�"�m��������>L��O�>7 ���u�2��Л$��&�$�g�蟼��Z�s��k>�8P�e����C�縥"CC0���lWn� �\������#^(�sD8M���{�߇\;կ-r� ��2r�aV���d�A���TR���r茔P����6�|km��I���w3��4dx>�&_,��{� �&���p��iv�"�
�]N��9�����nG7`T��-xQT�m0�晇���	�h��k��J��j��������dQB�����/����N�s�����ŧR����!!{�E��Ă�<A0{B�|�#Ӛ'J�AM���B\a�!�/
���Q�]at��z�VM���t~xi��>��������`<����+��跑�h<	��E��K�^?���n�R1�4:�.�5�µ��A��)Ӗߓe�D���a@Q\*���?�KJ�Q�b���-k쫵Iy�C��헄�z7�z�</:b����d�wf��b�uW�Sf#3� ��Ƶ�+�Q�q�ޕ�d����]�moi�D�-	��?�w�Ps��<��m�'��e|Mڗ�s�ޠ���V6������YuS�3�h�ֺ�V��*���}�PK�4zd���_�~v�^�>0;�cĈ�$f���k� �)Z�nt4���C5Z/$۶s�o$3Ix��������þ�Q	wY٨R�EE��2��*u���(�Q��dۃ �v��̲��9���e���nZL.d=�k�x��zv�^}�/������G����y)��)�G�|Ē��ڟ�j�@�����o��ۯ�Ұm�H˚{r�:j���y�3�}j�ve�A����<�?���t|�]���[[���A�"���:�p�7�>�R�/Z��%F����Q<S�c\�W14�V��������P�"�hm0j�����ˇ*1>D2|��˳M�����F�"����KoP�ڑ��*_�0��E�Ȓ�[�>��4�9*���;��:4� G�?hk��Mw_�O�u�V��M�ײ����1N������*���6���N�ͱ�\��|]�U���ȦOs`��Q��_���m[�I��3� =�˶ہ���,~fLJme5�-��C�4*��ӏa����/��2�v�s�,�o]�z|��}�-Y���v|8?X{�^n�]��DTo�r��,��x|2���
�3y�Z4�B1 �Q<FK����#���ݖ�c*Zj1��kq���<Is+���Ϫ[�F�=E���p�8 �?�G@?���;x�ӭZMI�/h?.�Z�̵�4�ǕV��J�����XM�C���VF�8��`�I#��^&�Y&y�4FFϤ	<+���,��<�x:9���<�?�nPA�0�6����v2ߴ`�J!��&��b���o�33A̠@ԉ6��:ˉ����KgXI�A��/�G!����F���~�!~����|6Ӷ���f^�w��z���b}�0�O̫B�����7�W���z't� '-L��_��n֔o��>�h	ρ���f5�y�d��BrgN�{�C�0����W��Զ}�U�P�ر�������R���ӥ��G��̰���5Me\)��j�'V����Z���b��#�c^s���6��-'Yʳ~�z����������!�ҞF�dЏ%�D�Mvρ�_�&�4�e>���PVQ�b�8�b8�HJ&i8	����R�'�U�΋`��{^��ɷ�#�����)�ƣv�()�]�/��A����Q�	"��o�.��K��u�Bt �����U=l=N��@@�{�V;Υ �<RJC�Jjߦ�Nu)~El̠y;)hWH�e�Y0��=� Vp��;��]q�:�c7�h~9�oA��`��W���
v������o� ��Mw@a��ߛ�v�^�����S�6�3�&ZUj�_��nl�K#ٖ!�E?f����JeH��m1Kd1Ec��N�ϟ�0ǹ�2�f�0 �����z���G�&"���]l	WY8gf��5�΂s���&���]4���7 4F�)Ȗ�k/�nob-�5����<�AG>f��D�b�9��	��ñ�;�\{Y}�0�6�̝1�o����S�1��P�'�X��^�m�j�i��*���(͈��5D̬��Y��W@�! j�4����Z�.���G>|m�H3��mn�C�3
�ZJ�	om �F�4���<�<��2Wp<�F�����Փq���i/�������~�=�����n����]$X�s5���=&���[�VD����xj_�P�������'!</����10&�,��h{��]"0��*:���,�ʓ]��v������iǮ�;��bC\}���+ާs@r�5����f�^(0,����l%^y^�2���`j|��*���~S�[��z�Ӝ�����jMs�*U;�\}0F���!Ў�Q��t����3-+$���Pqd��0��.��mǀ��� tL�ns�|3�Xd�3�z�=�2�p;�2�lKf����#���R#�2�y�tx��0T(ecf��ɝpW�z9����Oǰ�ףQ��3�y�DTQ�NK�}����NR2�����xUG!/P������~^��UOI��o��~c (R�(R{S�����c����X�#�.�̍@�s٧;��Ζ`�A��o:�-K�H�X�x.�)9h�W���-javi*�)�1��J8�E��r��M`�Λ��=b��<���|���BЀ�dg�*x�9J7�3��uM�Fѓ9�,W1B�4I2��qDA�i)Y�5I��ͺ���ฉ����_�%/��'��)j#��W(BZy$�s���m�^�>ϑ��x߱~{�A���9��@����V��"��x���P9jj�{F0�1�U� ��)L�ڻ��p��`�A %k�3�ݺ`ђ=��r˩��/ic~r���Fu����c�p�:{�.�h�3� ��^mܗʱ3�����@շ9C�E�Δ7�Jڀ��(����GD��=d�1�¾L���*��A������i��C��"!�N�] ��J����B�]��skR�yz��6'<P������0Ij�ԋ�c�ۡ�9�����4�@��uѼ5��=6�&�Hu\-M*�w��H�Ұ"/�BD�!=�}I�m�3{0zM�Eە;[��È7N���!�E���5�j��O��x�$��� �@Z��w�'�y /@��'�(u$�0�þx�c���C3{(�4���d��υ�p�}��J�-��da��4Ö�y�)��v�%A��A>HF맏E��D�f����{�r��Y��{f^�B`~��/����bW��y?�W���������d����<���R�;5���e� �V�=Ug>���ʗ�K�=1D^�c�(w{Z��������C8�U21�liP��$K^RI@�Ͳ�~_���{`i�8C�(?