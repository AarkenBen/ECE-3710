XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z~Oe䤗I)ņ�dә���R��H�䦌u�Y��.�S��w�b��芋�-����4ӵ�qݖ��7�9l� LD2�O��p_8��)HDg:?�adpU�!�w�+N,�Sdo+Lq[�}}s^pbp�ȥ�L������y����?��v܈���$'��J���X �s��B��[c�#rf�q �\�,�J�O��]Ҙ/�E3w,P�Ҩ�[�1LL�Z���XYkv<-c��N���q	D�W��g�2#��HG�K���>��)��g��@36�f	)� �f���Y�$�W�4v��'tW�������r<�ҹk#b������(��qA�T\�G*D(C���Qq��Sn)��BGd<$��C5���6L��]����xϧ@n�SdT�{=��l�Ό6E\=
��4�'���_�r3[�����m�E?*��LH���)�J��e,*/��9�Q�=�<EE[С�$��=���C��ж^F]ZH��x�D#/�!�x� ���Ѫ�C�	q`5	�~IƗ�l����<����x��a�b�GM}ֵ�вH, � �)�^�:a11������7ݺ��H�V� ����Ħ���ݤ^��[�]������a4��#S�6������0���i�vWcӮ�Z��qܝ{N���ID��dj�^���R�����Jqs�7�������`=a�n=f�UH�SB�?�^�8	�P	��c{o�u�-�	����  �yE0M�? ����#XlxVHYEB    3042     c80{�&��v�$֢�M��^T<㑘־��̩�4"�X�_V��'B�1`,�y�PI��F#�NUΦ󡑙�Lw�W�d����w������= �9$~[9f�a�V���Ϻ��b�tJw�68�TA���vT��^ǈ8�|V�2�r�4.�֠�m�2����@��&�����w	�c�u�"2(�>J%�$''E��3���lbGtOY��f�_���Hi���g����]�R�J��v&��?�J���ǝ���FLu�o��>:�of4_�!�~<!�확Q��
X�;��y�2<���3p+�xf1��_m�'^��<�xp�;0�1��3�]�'杩�ّ'���̀�}�`�W�u��0V�Eg�|��E��S���%���dπ��>�Ȭ]aE��4����L����)�T�!	 .���#xA�>�$?%�$�	V0�pJ�����zx���I�9!��Q�T�TLtO�ΐ�cM�����5���55��@_���n@�pߡ��eڬ��~Uٽ�^�0�G��;���HL�^+�����)!��n�[�gx9��M��8�"�+��ӂ%�JX���(�/g�%�5�k�nq���g��m��Ђ�X����x���pl�}ýT����n)$�E��ʴ�6���=���0�0�钏��s�3hC[_m~�~'��$A�**U�9F
�����)T>��ˀ�h�L;���GB��!���S�(~H������{�?�Ay���7խq��;(~��RUwd#�I���e��DEw�k��'Nc.ԬȪ��,<��&(6v��?�C��D���I�vj��7/�m��Z�hr)�Gf� �c�^]� ����9���	kA\�2�MH�R�1I��KP��Y%^䖦�W_�����#C��������Ei�,�g$��x��ԍ�C�%�{W��G�+��d��LЖ����È��f];���'`f� ��4��@�Џ�_kԂ���Z�T�������,��v�bC�
��@��5s�ܷ΍����>�6��94�:�0���ظR�����߃�9���*�"���+U(�4='�u��������y�G�]��&	��!�f䆮mV�l���o�)��L����c�ߤ��0T�6Eb~vI�Ja�@�2}ݡ$���������B�ꭵ挮��!pA�h;���f�q�^9/G���p}SZ��yu"����	��~2�ʲE�s�&�m�)��CӶ��7�y\����T��6JR�EF 3�O?j��{~./rӨ)[!��J�e�#:=���2�+��@rf�9�ή$�1�0�W���M�ٟX) �E�ǽ-_����_k	�(�S�W�z�)�2Rf�ܻ|b[<���߆G����I{���Z�W/-���(s�?7�7ͧ�h?�:[�̱ϻ{7Uh���s����u���1�cN�Zi�y��l�x����A��&u�� 
A�d��:�Db]�on,t��b��$���Vi�vkVs�����0�ȡA\��_'���B�>�|��5[���6��K���������Z1��$R	u�d�)΃cM�s�-��]�Z����F��mߎF����߭��E�~�=_�ϔ�H�3IY�)V��4*4�N�SgT/�5�I�El�}g�ؑM�ɴuR%�[���x47���t̎�4n�/�&��5T�x��cwt9�4�}!O���7�?�B���+�.	P�3<�2 "����sp��E�E'�u��F�"[�����ͭ��-�.��Fp�I��=;W�Cv�@Q�k�����Ṩ/�y��A�oN�X�� �����ZN�}��h�dWu���!�-}$��^������X�WW�Jϊ���[
FGy2|p�I�w���ap���p�*ˇ�s��7��|+�*�L�a�,8��JX�&��L2� �B��Gb�"�ⴂ90TM�2�Ɇ���
���I�Re���N 3×���9�m빮Y�0ܡ�<�>L��>�V�p���a��b7R�?![��lBַ!�q)gS6r�� 5���Q׷�`cK�aHLü���&#6U%�������#8� ��&�"��QӖ��G�28��K�]b�Β�"�Pr}������b�`�����,�k_3nwͺ4�^�2��Y,>�&K�lt��_`:o{b�U��0P�I��3G��VnM�NQ��$u�F���\ۍ(�\�)-�F!�]�fQ�O��r�{��l`�aS<7'�P��JF�W�K@���р^W�=���]��>4�wh����S��0'np��~J"M㈶�m��s�0�6��ˢk6��	]�
�M$�=a�Sgۘ�T��/n�{�o���2,Ӗ��H��(zٌ�	�Ay�0��"����kZ��۫��Ì��]�!l i���v�$���N��۲�qA���^>�G#�h�37��dU`��6u,�*4\�E��P%��/��0Q9���g�M4:辈h���m߮�cº�	5���O�R$c0�:���~b�#��VKU�>���X���E�Ԛ�KN�
��`�=�Y�e�7KQIK֥r�~I|�Ѝ��<����,:=��.z�x{kD`g�)Z�� -�PhU��Wp�a��R�,����X͇a��9��:-��H�p���R�#Š�w�zU:ح'���{�p���p_�տUsu���L������@�'aZ\�`�5���@Ƭ9���"<�2�����c�B��&�~��j�@�6ȩ��W�P��^5m����)�a�uBN��/���h���O���Ȇ˴	`&*�����&����	�jXw�1��gj����i�c��E����f��;���n[P"4�7i�}X�i�~���,ef?��S:ito�Hw�D�]��[-]�胣����y�K��w��yv��B��<�����_F�!�F=��:؁@~|e%m&�H��D5ba��2���Vז����2��l/���BM|�qݨK��Zwb��)\�˱����Y���.��A�� h���\����J1�?ŰK	gn	 !�����ŰIw�I-�������K�֌���E��P �$�[ѥ�,, z�Ԁu$�le���t)G�ޘ[IĨ��N�����,Ӗ���sW�V�Y�5�i����P"�[��J��JL�S��e�