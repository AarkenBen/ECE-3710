XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���g`��e����_�R�f;�wȷȎ�ոD��wbj��}+ef��t�R�מC�",>�Ҷ�.[Hpn�]���=�����=Dk��L�䲻��UHY÷Y)ڟ%��C/�d	O�� ~�
�l��V��72D�0.��%��6+�8ě���{\"����2����l(��=��!F:�Y���N�] s73��%����x��ǘOq�����
r�}��\��f4}-�0g=R�~�7�������A��cli�c�G����m(�t��활1NsQ%8km(��p�Ǎ�\��Hh�ZK����ѲZ�um��,<Pk�-�^�a�DLfVs?
�	8q�}d�b���+�
�׹*-�#߅� cèn��E����U��8�z��	.�\��B>=�5��Y�S�?�����~����{8��ʑL*��wI��F܂��:��8��+e��R�o�� �*�GP��2�bž��Ά��o;o|��Xl�kV>%1#��v�9
��:ZP����:�H�M�ޱ���"�_9��G�q�3��z����Q���!� ���6UvЁİ4߸ ��_泂_��Pd{S��a.F�������#w捸�у���TH���C���>E�g8���1�.�5���ĝ�K�3y��C��y��J
�_
�'�aAM856��s�ـsۺ�tv��R��9�"��c����ֆmEx�,�v��r�&��Pc�.��4O�?=)����K5H�x�D�P9T)�O��8á�uti�|��~�XlxVHYEB    aa31    1e40nKd��t����'1U
a�Ȫ�
��d�$8�8({�����~��1�Ro7h+d��-��R?��C<C�.Z`x#W�q��,8_���G��FǢ65��Q+ʽVݗ�Ⳡ�I�x	�V���u�>p�ca�:��6m �O����1�V�|��Jv'"%���&���nC)�3ȈJ�a=D�n8���яd�@a�r�1�.8>f"a�01��A�V�m���o[g\\A<)³�j�@A�&��%�q�%��,(�}�������}#?�-r "�?."���^��z&�H�p���,�;�T��
g$ϻ�dL;h�Md��P JO���&mRBNt�vϚ�RS��)�3�b u��9���>�ft^C���	5�L�Vz3����Hդ9�[��r+���_$��վXF�1\��$Z�E@�%d��"^Y����$��¬�(S�x<�MH��-X��tV�����a �����	A��S&*_�jt�o���ɚw!I����f�8���,�i��?��~���
<Ҿ7��V��<'�&�mM~�1�i��A�S�����.�AOJB%��a��E������&����H�5�!����^yȿ���)�&�?�=1@vg�^�O����˨E�:`I<�c��عjO��U�V y�k��K[�X>�urW ���ө:��-�^nݷ
��Ud��n�caB�:+]:�5�Rc����;�#����//�>@�`N�I��AP"E�c�}E�p��: g�3!���)�����ʓ�iM�g,�:���е�B�)/�a9ڹÃe��@6d����'F��"�����>X�od��8oq�S�A��� k�����kB1��<Q}Ll�� � ~�i[幓)���t��PTl ��^��\�����k�:�y �o���3U�_��{WԴ5�X����\F9�G߆�Ν�w���6���¦-�K���y�><J��l���Z�nb��Tٰ�L��
H�"�N�.����Z�u���h�6�kI%qh-���I�η�%A"�Է�=�[*FZ��0�005&�M�=s#����o��3�<50����/��b>�n_���@���a��3c�)����|�O�o��S��$To�BV����Ȱb ��V���t߷7��Q�[��6��ࢥC�K��m�-4?@L��ӣs���"�Ǔ%�@��9P<Q��~�
��`�iZ��Q�{ ^��H�v�l$-� ߁�.��>۫t�SA�|����w����k
<��u<���IG��h������k�/�7An��7'V!�l�� n�7ai�������#k���M%� h=��P�P�x*u��{���ZC1���}�.��K�,S!G��A�"x��̢z	h�|���B(ص�ң ��Xt[�k��%j�G݁ybW�u�e���)��4j�R�E���N�%Qd˕���}U��Sʹĥ�;���s6P�y�.J\pF[��h-�=�&d���5��S"�Y��-S"!��/���U��b:@V|�ل랝��X/�҇�<����g���{����H�S6|�IA��cE�`&9����/�����7zy�(7�賲Jغ�\}Y:�{`0�Z� �C�!���<�Y� �<S}�z��.ڨ�����	Ǽ�~�֜�m�3�;��帴YW��~�5��*q�����U��	�r5?���(m�s�n�0J�A�
h��7�G
��U�j)�U�1�y�|��8�:��/&<��yPǡ��@�ߖ7ڨxzѰ�G��[��^-��.ֻ�(6��D>eʤ*�4�f��橄kl(�e]i�&�)��c�L�fe��
+ fZ����!�P�2/�?����>W�k`c.0����8b�7vC���C/�ú��"?�
���fs�������h���O��l�]��	!��U�fp�W��>s��[���o�E���>1�E�<�*;_S���0����p;��p٠��$��^���%�h8yx���1����}�I�Tv��i�w�SC@�n#����*n3x�%⎱Ɍ���,te�M�ʒ��x<�|2�֌k:�C6����1��e�"H�19���_��k�uI�K9]��"A@�'b����7���\A��<�KZ��O�ě*칡��&�_ ���Y��M�YW(]���J����p���9��0���R¸�0;����nW��R�{'P_�1Z"^$�,�5�gl�ǎ���U�w���	mE��,}�\vF�ᶑkI17�?e8XRQ�Q_E�ǔ��.[&k)���ߟ�/w���yL�}f¤���������gX5�<*iO�����-{
'��v 	o|2N�&-~� 5U�v⁹���E� ؋���-M��y���#.>j�'ט�-�|N�����./���]������'
(�6��U6����K��޿���(��*S>xsQ��i+�,���������*��
[�Ŀ.�M��������U�nji��a$�7��a��u�Sa���:k����%��Q��}OO|׻���~��OZ��WӜэ!�;�~�Rwz��t�n8u<�	h�]�o�6�a��ӱ^P�/��(#OQw	��<~�b�ņ-9��i&�V�bz�]����xJ��ݛ�xĻ���e�z�qi��?Qt #��� ����ۅ;����ꕌ�"n�ny�gS <*�5�J`l�r�x����m2!7+��'�$82rf�8��\;�Ăa�SZ�[��5���w�I�{���Ȃ�~�;z%BRS1]p���tٴ�Q�n���jV�a���J�pp W�K�n[[A�D�40E���}Q*v�}��cp�H~V����Y��,�k#Yu̴nKnj���D(-c�5��h���u�,�t�AӑH"���`zԿ��>M�$���l�q��_�:s�mc�"A2$U:��I}R���h�dJ�,�.��5��)�&]����I�'�<%w�e~�ã��eK�_���a��C�j���l��E�H��|�V̇�y���F*�����L�Cl�-����q'��{C�=�ރZ���bƁ��Y'eA����# ��E���X}F��D��.ӎ�L��$Ls�X�X�ɗ�'�5s�\os=y�L�˕hvf�t�E��@1~� �G�����Mz,�����ME�#Ҙai�%A�뾀G&����QG+D�d�q�.��lA�� )`ߤY)�nC��+G$̇y՘a�vLZ��f�	��� ǐ���mg�0I��Ue�`���^�J"(�*��l�(�J
Oh�>Mۢ�d�x{��9a`#k*r��j�>�/ܘJ\��#�U���!4�L��Y��QGg�����,}�B>r})�����yH��ac�%�nO�+/]��I�;�egx�+>,�#`��1iPJf��_��z�l�޶⺆�{���2�049�I:��F�K�=���
��a�4	���V�O�k������a�iC�ŀ	ǐj40�i�?H�<2:I�U�lTy�	9z ܾ�ú�������[b�ݪa�>j��H:`N�e�X�(27�n��F���l=���#?%�o[J�%�l�W��Pڜ�|c�a�tU���f߶Wk=p���)x��0]�ǦN���a��6c*cO���R�wS���1Ą�Y�?ٮ��o�����J�K\ܡ[NT8��x�b����6�P^��3��կ^[��-%����s�h�c��Qʊ����K�͵� ��R�8�A�P� �L�c���I�U�&R�� �2��:�\�����)�zռ���5W㡆'��z����M#��(�Δ*q8w������E��MK�-�7<�/51�H`��+C�eF�MZ���ϗ�Oh���i�}WL�u��W�,B�	��
�NᎣ�R��S���=]�63�n-��޹�=y�g�#H�7��k_�73�����͟��b�����4h+o�M^�4XU�6Q	A�F��M�"}hLM :'�U~=�I�~�1)�NXh�F���]¼�������곸�_�P�������%����!�a���AI,�Z�:C*� �Ƹ��V|��[M�!���]�G0��/�
;Ud6_:�V< |�z[.����M�|k��>�XrX:R��y#������'�o�F? �Wk����/��ˍ��"O�Ը�\�?�ʇOҰY�C`|�o��+NJK=���C��V�׬�Cԭ��P�󻀓.6E�HҮ��%~:w�r�i.���,��g�Ğ�3���A�S7�<�*S�Q^
��6�!b.�+O��!f��i� #�W�YkK2s�\��Q%+���^��h�Ӊ�D��ĸ��Q����g�p�c`�L�SU�O����=],��* ����.IqQ
C����]����?J��ݹ�J��KH�.���t�[M�q�p�	�7���V�� ���ut;��̽欀ܧg��.e�,D_�.Y�"����(����$z��?������"]�C�_�>5�xZ!��i�������2��E�4��7U�����o�O�ყ���B�6*�q� ��;ڧao�e�2�>EO�0���|�,���z����Jp
V���\���;�@}w��D�7K�]!t-0;]}�c����ܷ�a���H4+M1�_/�QL���7��A��H���N��-��Ȫ��XFl�q�%��>Aͭ-�a	����wXҢc�C��'xլIBv:��[T):SI�p'=�(f���]"���*�Fǭ�O64�!x����o��z[w)ݿ'3���C2�=�{WZ�'�{a�i��EE��r��,Q�X'��d$����;[r�BT}���*¢_���zg �E�V?x_���ivp��~�m${�li��@����~~rw��V��F�����#�x��e�����Z�#'z��Q9����,_���%mi]gӤ�M"��R�l_ӳC�u�j�*`m)O�x���#v�Yv�J�-hެ��9�=̡�����^����]Y6ˆ�"'U�Zw�>�F荥L��k����r��Әɿ�+'���+��ޣt@�ZRCt
E�l�܈��J�+:�{$���ùe�;#縚k���?�R���56v����i���5��ɟr�^9d�W)��3ȅb@�L���2{Az�p?�А�#g!6s���W��\��5�+��fV945�[a�|	
2'��qGBs�X6���������X]9�����35���}��X$Ԟ�D�k	/e'v��ARŢ�LQkM���L��S��:�3�U>G}� e�{K)ZR�[ٸ\C����8���F���l�EjY�E��`�����!��
NhJmV\���暡�$w��OW�uA���͜�?}U��%�7�)Q\y��{��������3����b���)V��u:���Q�#��m�m��A��GѮ%hdtՅYY�9l-�ͽx1����n�a�ȗ�X��W�����$8�E�t���Az+���k���f�J)��D�1P5%��YBʋ�H'�qr�FH*�F*�7�tҜ��x�'V�b	���`��I���[8����;Y�yK��꒙Le�ېPbKh"��Lf#�8�;�(4�Tb����8��snu˴��i�8I4��s/^L�v����I�ĺ"��zS�+w,'_�3`��Z�Z* ݄�1�o(�:�/__=�iQ!�%�4!�����#q�m"ηp9�|��U9��D�
�~��R&�Ϻ�����+S�_�栖��`�YDa9�s��g����(lh����g�%���ǥk��Gϴx7=�Yk���ù7�2��B�@�?p��,����,�`4E�g�\ce�	Kmn{��qC�w� ��BQ�n��D��Ý��a�����)¨�6r<��� ��B��;� ��2�0��f&�@�l���^���m�m�߽X��`;�S�ل��v���+Q�T���>˯7ʄ�O��|,
�����ǋ���b;ǼQ�u�(�7�ϳ9HHw�03J�(���@.ɱ3�������w�J�՟�v쑜�!Cp};�x�!"������hx�k�৽q�:`K`Fvϻ��Ĕn�i **�vd�7�k, P�1�F�8B�zS�~��^�y�������U)�'N�sĦ�L�"[,�EKo�Ćܞ
\��Q�~+�T�r�}�om.&Q����+�p��N'�޸��Rf�����-cd�lC}���.�!)kIkn�_�G�lwQ-ĝ�:쏷�K'�����(�#���al�_S��33�re���Z$����_��]` R�	Q8g���K�Y���x�Y!�)'k�d�D�'���#x���]C!�*J�l:�3LB�O����)�s���M�qq�h�	�.�^3� �H�o4kϠ�Rd�f����+����Gf��Ќ��2�y�Y-xB'����$(��;d�h"t<��	���A�a ���LM> bBˀ}�@�9Jl~�dOg���\��])�y<�^�b K�eD7?�{�6^	$Y},�v4�쉪�M�Vn׼-!�2��M9>���ߋ~�A�,����;�N�y\��F�m^86�B�m;�_g8:EN3a�Z�A�! ���Zߒ��܌OH��2�Ō�yz7?�ǲK��9��Rge������1|l�v瓖@�0.�#� S��f1�+xXΚ�+��$�X��������8��j(V�+'�:����$�'j���s�tzl �3�Q����T�w��A�35x�D�_�I�����2��!K�^�݈�Tm:DO����,�|�o�~�v�~���ި�[l�x���2���v7�$p"��7��|�e�Ap���ǒ�㹶�)����o=dZ¾&{9�1��EԦ'�f|p̺E���
��-���s @k\M�>N�k���,T�d�E��*wn8/�vct� d	�J�+)U�l�|�JM� �Ԯ>��� �Ѧ��Au �S��xt�9;QCfw�_vp��[��8�у�z�)��`����x�*��	P�(���F/���@P�aTr{ѭ�y:24�d���N��Gom�1���p԰`�$�g�P|���i'�=X�Tt��V�p$��!�
�
 �s��,��I����u���N̜uTR��G~o��g	��FH5��I���Xc�1C�?>xxՋ�n�hSL.t;B��ϑ��%o9�OB!r�J<�������u?P�p��̞��x�0�������j@�-Ro٥z--�݆m�H�M�����=�����e�N��a��׿u��;���_%f�^?���y6�a_X�ܮ=��oě0i��pj���}I�P�P~��/Z)�:է ����#%��mZ�w�^/��3�01���bVgȹ��;Z�|�:c/�t��G�Q!�w�\-u�N;L�#X��v�X�����tt�Q���b�� M��#����~*w�� ��m�� ����JO
��a�uG�A?:?���D�O��CB���;� �����������/m�@lL�G�w�+�����߇�C���#&؞7G��r{��+�۔�M�]�j��'��R m�1UW�_��&t���<��s�\���Ԟ�K��E��g�a��,sc%:5hՑ,����o���*y,ĺ=�
��tt�ъ$�u�T�(A��f���.R��|�B�qьC�g���;Le��Ӕ�a��J�-�d����Q��嵹�y�]vp��k�{