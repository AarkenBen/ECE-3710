XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_݃�>^V��C����"܇l<��(w�EIM���?�k:���9>��^S5�H��s,e�ߊ�y�(�bpEw�Y����iP��t�ck��V��5 Uܘ�E��Xm�t�!��F_Dkp���4C#��6*w��6 \'|��}7�-���D6��-�U:}bڍj��m2Ŗ�J��ƫ(���;r�E�v�$b񛳥a�R7a}�o�O���םNF���q�A��ALl�I���;'�4��;�=i�t�s�r�<
��좒oϐ������;G�z���V_�D�w.Mu�|'�2����	�M�U}�;�M$�T����Ą̈́�����v��B{BI�^�3�������?+M�SQ�s�1LÓ)_�aZ����e�C����<�sG��!�l����GvK~� 0,���Q�w1b�)%�M ��s�رzњ腏a���Q�v�ɇ�H1C�,À��9�����r�)N%��3�]��Xd�i��1�U���۩���^[n�ġ�Y1*^�\�ul$dX���;e��i#�׾��S�z`�%�}b���Zr����Í:����:!b�4B{��P���~v=r�U�OvW<u	;�K�(��x,���nr[[��;p�����$�"��ICސ�l.3'Qsǭ6�g ���{�����~Si�y$�!�=Ϣ���ְ1{y<�Q��^�/�(RI:�'C��W��e茖�m�R�iQ�a��z�5���w"1��~��u��w������η��:XlxVHYEB    fa00    20306		��;!���b���/�9�>��3�!����``�"|��y��Z��7xp�����+b�n{%p�R�"��N��8]�X�a�t�k������]�r�%Tn27kr���تM����o`�V&�D�}9ѣ7K*�n��%���Q��n1͏��/e�mI\ 6l���9(������~�~�S���+MtoB#��b���3��-r5A|��
O��"j�.e�Y�אLڲ.��}����#���vE(ueI����C���v6��̄GQ�O�@͉�wH�֧�`8.����lg�*�ҭ�&h�*"�X3�s}E	4C�/��q^
܅A�m����I�|�|1n�|b۰��D=�~N�]��Ihجh���(c*�k��^ށ)$5��.�'-�7�W`���s~�k+��f�/�Yu)�W֯$g�I��7Ȱ�2,!��|-�ۛ���{�G3���׋㱜;�d�D7��*����b�>o� =V�f�9�`�	��% 2�#�`OވKx`�lw���Je�;��$��{G�}�E���C��B!��񨷐�3�t��ip��̅|�����2)®g���������𧵷�?���υ����+)�tW�h`pza��t/�E
�
`��T�m�LI
=��j.�Qs �{X���;s0��y{]�l7�;�IM��h@Fx�?�I�����1�$���輮wbD�&����XF����Ie�U�54�ozB�g~�H^:��s��M���w��h��6g��#�?zA(n�D���F���#�n�hr7�K{}�xe��;�O I�RN����gsJ�	�
��<��0ib�DW{��Q4*�y��5��[c�Ja0Mچ���D:XO:3&���Ӟ�{Neo$?�̏�70F�+��~���"�$��>��e�ڒ��	@Xݵ޸�C�۰�(��~5�'x{)��(��XAvT�A�#��S@KPf����HJҬ��I������e���j���W�?�sٰe��b�3��H[Ѭ���5(/���9d��z��?�&/�����#l��B�����b��7z�ْÒ\��e	)�
0C�C��U���g�]6e��XWT�Hц�r(�T�<}��U��-��Y�y��z,j�)
����˽Kqa�c�eX]C����e���3��D�'q��.�C�I�w�[zC� /���9�z�� T�x�ix�W�;z~����ظG��6G�Gĸs"���)�(��t�����p)�:��T�خ�[IC� /D�h�x[Ǹ �	X|K$�� �,J�gtm/_eF�$I
B�������l�����r���_M��?8�����(ޮ+�[���B�J��,#pL���*'�F@�MH8�W�C�ت�+O ���#ez�aO�?I�ET�,�<���9���@���C���`�7��<d��5���X��܈�#���/m�Ɇ1<R�������~ލ�C��4{��R�3|����1���E������ti�>Kɲ�.v����H�lFqi�M~��~C!��lEw�^&����/������?�䆟"
�_񛿀I�1(�D$�k_���__���Cx�g�>�F��|�k:k�%���1�Y�}Y���&}T㬕��+����m(�M(�O ݡ+�!�� �=�������oI���0wN2�3��1��K_Uh,!�@�km`8#2�������L���M2���>����^�9H�[� ��L3;�=�dde:Bm������|�j�U�I���Q,+�K�*b[��rR�M��� ��rO�I��-p�&��n���m��$0,�P�f��Z��ÿyi��D�ӛ��P|Kn��ˉ~*R����J�]Ӓm��|O��������%���U��z��o]TZD������n^�4�O�L@�(���\Fs2�9[�V��z�I��R�	�8�ܱ�����8��~���;�лK/�`��n����޲I��'��U&@���l�ݽK�/������ߑ^uZK*��/�>�b4��?�b�S��opַ㡕/W����%U�'�a�Je�<����r��4)�x�(�e��h�m��E�e�~�6�#�ZYtp������e��N��4و��X���Xa�R���������>�y�A���%�t�k�~��yˈZ��r'��`^�Jش��Бw�JP���ȇ��̸g"�����.��(�U�^��`P((7��f�W�Q3��wtIv�]�	4B 9�ڬ-�S���F�#n�*j�H# �(���Z&z�Ys�����rt5m�.y����<��;�3Zl8�\�p�J�Lb�֨���B��ol]Zܴ{k}%���2΅�.+1U�����x�����{v@}sZ��NZUW��ߠ<�ݙ����q�XG{���X���g�����q�+�q���`@���m:,2��]��Wi�Li������Ծ��7|����u]c|�bZ�C��-�^�b�ܖ��&�e��1@z�3�3Lmf����T�'���%�ڰM��T��v �a� �\&���6�>Ѹe��
t�b�S�f[���ť�ޭ�$����s��(h6���}���Z�i�W�]"XbKם�6YQA�@PwR��)&{Z7r1����7����y���0�C1��P%B��K5-q߂v�P�*K~�H��]�i�����	&�OZ��ˊ��X8�Y�՞�5���r/pT��?��&o��5�a%�B~���p����ع���%�r���A������@��1�>F�����AϜ���+��<�� �f�E̑��>ó8TM�̌[;�q�\���E8������=��3<��ʍ�����3od嗍U=�J��\���������F�����Sц�����r"+��F��f�89[9�|b^ve�E|P̟�~�h&��5X�[6yH��\�᝷�>��n��SM�Պ;�V�iVL���~W�Y�4	a�!-m�:9S]!�����B1����[�.'�3�;X���R?�����\�*�}�DtҘ:�#�S��lY�y���+{XCS����+�U��0���1g��3�:�QEE�K�o</2��.�%M:�?*��Y	Tx�'�Cw4�UR�[�	u�;���i�?Z��v!����d ��ء1��N��O	hr����'��	�/]�?x_�S�xh$�K����X�b	_8���H���whV���*��)G�H��CZf�{�W!?*p-eX6�$Z��h(O0Z��2@��}.��I�w��w��&�F��ͤ
�F0h�n�MW��vh�{NK���|�\�>�I!ќ��"���"j~E[�>}���yA�~l_q�7w��v���0uy���Gp%��=P+X��nc�=��=��c��Ip8�y�m�)��Ƚm^�(N��֛�.�k�[%P]��0\�<�=��b	�-US\�8�Ss#>�f���*:�q�*���r�����'g����$`fѲe�Ǉ|�Z2��r����><,dfů�w�*���ř@�����Ltk&bIإ^�`c�
?�i.V����<��b%��&�Ḙ0[\��*G�x]2��$AXL��=��v��H�P	ӓ(�I$�<Qm���x�x�ʪ��@�}��{x��.���mY<��-�]�ؒ�:��$��U��x�Ke����ïH��?/[iz�Y��N[�-UNG�U�TS*�'~xX��T'��ᚊ.��X��}[��
�����T@h�ӏ�O��$ReI4��\oK��T_�]��$�ì�'���*7��#����m�?���IKEH�Kk��W(��S,��
���v�_��+X,���Yі�d��T��d��@�?��}m�������#��c4�����#�5xWM�}�.D���4s�q��d�ڇ�4�����*	��P�/��}8,ٝ0��0O����7�,�2!X3&�.��wAxb���|4n�tۀ��4���5%�/�ͅ�Z�f�E:��!>����P���?���4_qϸl{P-I�V�MTqi�*�&�.�C�C�n><DT�zA��(hu�[�8±���O�}�<���O������	xp�$CR�\�1�\:��=����!�t��1h�48hm��1�l���h�{!?[+!ɹ�S��Dڄ�|W/�'�X �pz�<��dH��wJ8|:N%F��@�I[�,����"'C�/Md`%��W�?��px2]�${$��v�&9��6ѩo`#�,7I6��h��e�c�LF��l����|Ξ�=4m���f#c���9�ݪ�O�2V�ֶ�1j��/�_l��m�:�P�;<�K��y�X#�Z@�b�/���T0C|/�eUH� �My�H�?��,(����_d�zh鷪 �T�����xWr�mO��OQ6�_�9,pe�0�F�9���ʴ�K>=�k�C�ST3�\
)Oa��U�P�e�m��x���5I�)�d�/�xbUBV�$�[_�;��whR�Ix��ײ���u�%���Y? )\�E�����=�5���W	œ��+���S!�2=�U7�51�I�p9Yn��zA>��I��eXZ��� 1Ó�[Cy�R�d�N�����,e�>�Q���k���!`j���h�܌�,;���G�5�:6m�v]�X�Y���2# Q��W�弌#*4��&p�ev�t��ǘ��cK�Z&�|`�By񭷷�%��1ɔ�v�D,ۜ���*y��^���`��Ul̄)KWF`�v.��ͤt�B�vw5�=��X��]���hX��҉�tq\ސ����<�e��繹̄i��7Z�oǵ�]���I@�;ID���n&�c b�z�s���_��6�o����{��;O��}�U��>�3A���I_6ұŚ[Sq�M�u`Ŀ��=pQ���й�����s�s�j���}?�UX�ţ��X"��O��ub����?ֱ�D���E��Z�/�w4?�݈��z]H���kD�6'tûW��� ��b�c���@z[̄I�z���?(1ư�tu�<��x.�YK��8)U'8;�Q9&����z&: �(���p�u�w����j�-j%���T���nFY�J�
x�A���+iW֢sq:�m�&Ǭ'?�1s��yu@�㌻�t�kve�EVi�"��02�;�3Ö���*�J���`)��	�̕��qen_b��eeQ_�4�f�r� ��.T��S򏹱;��$�_X/ ��g.�$���v��)mŌ����V�bɜ�@0E�n�De�8��y���{>)�,Rd�.�R亁cEC�1o���^���F�����J/�f�VL��Tg%�v��ifhĥ$nDU�P����͞�`�Nr[�sZ۟�G,Ғv��w%;��Lƶ��^��ugOL5˥���;yLnS�)m�\�.�3�������s�ܬ�L�W9f�8���� wsOR�-#XsH����_ɉ}$E����W�7��)�N��
P녢�v�	�>�r 屝~�ɣdn���2GQ[A.��?ne�F�x�&�(��(X��% l�e��s����wy��p�̦n)���S�v�T��C��d��������qh� ᘨ���s`^�)�(�dR9T<���7IX��z���[@���"})'i����+ι�˼��byq�	Z���X��z�P�#��'h�>���DnR��]�g༇�� D�j��D!Cħ乡�3�5�����$�� _�*D@�|P���9��m�ͣ_,-�P�%��qX`�
:Tn %����;��� L�#-�K%Y創�RU�K���Pk ��@��>�)�����^�|÷���Q˯:"1(�"u,���.GSgb��_������߭c��>)Q�rj�nٜx�5�����/%�,�Ŋ5%�����d�RS���N[,cjno�Ӡ-��t�ݹ'��G�3"��c��@�g5¥����͸��3����g�K�>/�E��P�C	�JPC5^��\��!��\҇=f	$�Z�u�+lF^bٵI�D���aU���&���9f�s�ha�@���_��.e�ݧ���'^����O�Q���N�;�b𹊭���Ѫ�.���E�
�YN6Ź7������
��W�������P}2{�_�z�� �6C��@��L���o���:��qW���95V�9�!�h����&1���;��*
���'��B�{ׇFŕ�Fd�R�{��@���R>/N�q}����@q�?�P�6�	�c3��=L��D�tJC��P�޹#K� ��|VR���Ba��JwU��3�:��/��3s(؏Ut���גЄ0�7>�"c�B�Cq�I\DK�������Lf���� �=��k��G�n���=�{λHK��������Ya�s$��J<w�;�	<���A�"�r�*�T~b���g2�o��b?&������{m�����'()�c�����I�����WKq��OD';BEZT���$i�>\���CTiV��ݩ`_s����m������o��\��wP�4���2'1m��a�t�n?aF�c���>\�_B�}��R��#%�53{��H�@2ro��,*��f�(��r�oa�D�\�pA���r��͉;����	riB]�v����Nņ���ݮ�?�h�|�汌mE�@�'l[�UPC��N	a�� lL!];;�o���Tr�+_'On��Z����j�}�M7����a�\t���Ty�I��OD���jo�����PؾJ�8YҶ
r@/�2�~�Yq��3��Mݯ��	��1t�跎�:�MR�nw��ʼ�R���)�����
�>�M@�b�@����l��n_��I�ѓ:���n�<C�N�j�{
'��H:���}�[� ���@S�.�Vr&iFt��D	�U%�&��i�c@U�M3k�*���>��H�.�U�+.�N�|�02^t<l��g,��9@B�eN.�޳H�|�X`v^��-jɡ�\l鲕�lׇ�ȥG��@.f����.U� ��Rm�-��J��=A�
�����h���nje�[��2~���K�Z[�ޢ�R�Rs�2H�L�`��_�R����Ny&B.��mZC�î}7�.�(R�� �)P� ��6
����0�_ �e�y����~VxRzO3���됿��Y,��ݬ������\�*�����q�\�����5�G{�I����q�U�j�wW>��} S�˰�s�H_A!m%X$;�>����!���Ѩd�?��ut��M�^q}����3�s�E��m`ߥ���-�z�o��{aS�8��XK��钑��(��	p[���I�`�B|��ޕ�������b�>��� ���F�H�� �K SbDE�>���׽���&��5���X�c9+�	一*�$��
�T����Oh@��ꖬ����0��4�C��,�K�(��Tm�E�6��}��ݠ���~`bu}��1{3�ֱ��w,֏�YAO(�z`��BY�d?֏�+Y�}kGa�x׽������hp-��f���)����>]ܦNȄG��e����ʊ,�N�
�U��K,O1��c��؋�;��e]��J �i)˨*���5�p��u7Fm���L�2C����	zQf����t�{)�������Q��է E��ד�KL�t�Z� w*�~�"[�te���!�fCB�(�F'�GԋNb�e�g�`��ť�θ*�"y%dN.N6�x�F���y[���j��[��BT��(H��`�V���~
��4mJ)9~�5S�m�����-����Ð3ҔA���$�[Gk<���?�wZ۽�q4�D�D`=�!�#��3�f�V�\�m��Ms��:s�+�gsZ�~n���r�N��U��zg^�-ē�O�}�SV.�#�c[�H~]F�OMF��u�<r"�&w�(�w��B�=ϸ0ׂFI�^~g�a"��q���|$A3���:�&���bX�2�����KO�n�q�L*�m`࿋U���շ~-�5��<��凵�y�@�-Y1^[؀����Z��6����,R,�ӎA�j���&�)3c�>��Ά(2�i��l�(ts\��,��'�z	&P��Pձ߿B���	��SXlxVHYEB    9620     d70�e�X���D)o��`�
~��7C*�Յr[lX��zs��8��z�u��`Lh���]U���~K�fv�a���'y��"[�_Tre��m�C�dܲ�c��x����K�Q��U.cҽDK�pc���@W&Mdü�+E7�`���'�y;�x^lMĂc}V�GiO�V]Ʒ����O*'���i�W��Н�Χ˅���ob�G��#]Ita$l+�v��cWG\�7��Pd�D����!X~{,"�U�1	(����8M��я@���. Y*�m�~ɊUn�!�v��`��X��-� 
�4��*��b��19��p;_hZ���{=:�ЁD�r����K0r��]���c0��%�7$����+j���(1�M�p�f,��3|j
���f��[o�>6�O%M�v&�>�s+
�d������)��}׌OS�)a�-�>��U�u"A.#���o,�pr���ʥ���pX��SpP!3����t��!�s^I@�nC��H[��&(u�M+Y���oZ��A&�����	j6�섹�>�B.�hw����j-0�{�U�ym������>��i�'��!eL��ޞ!��|��-
�f~r^�c�f<bzVNtܮ�����/q���HuV����*"��zY�>~�V��l#�)I@7�yt���/*2�U���9�9x8��!_8��F��FK�!�;����X���l��w��8�0 ���s���B��P�K|���͔��Qn�4s)�qQ�J��q�9�W�q���F�(�b�������+�0�s�!�g/z�;9"a�j0$��Cr<H���v�9w�rmݫ��;B�x
0��_�����Xe�h��_G�d�s[9�3 �L`����A�)unNF���5��r�F���a�ߗZt�����2g�#���h�1�92 K��j�Q�r�sG�+
v�b@P�|_WD��2�s�+7۫���3�
�kW�@�=��iJk��9�-��g��6@�vw�	�X'��+�v#縤
\x=�S:�'0t��B�{,�� B?k�`���� 
yxd��3��Qߪ�� �g9л��Q���^6�"�sH�4e���BE�P�;L���*6���]�Q/� 	)�(�]99U?BR�7ۘ�|S�夨���)�C�bi�2I{��~�y�{��x�h��4��#l��K�H�>��؝ &6�[]��hM���	�B�{��}W�b����%��-Т)�T�Fi����k�/� %���<����IU�Z������Ձ�"H�d5�U9k^��p��*��k�ޟ�ra����te۬�-'�#�8u��h��'���+/do�)V��'7s�Ļ�q���I����ԴT)�j-�շ��0_}uD]8V�R�?EP0h!T�U`~����Mj<8�Zq���wŅ�̃hO�>���-�4&X!�����������=V}���s�ː�{���@fRk-�u�Ĕ
.�pb�
�������`׬߄~�z�Ql������ǀ	'���Un3̖�D��:��'��ݜ6��6�M��N��'����74�}F��Z:�'�.�$�(3�_���}Q)�Q��1S��}��{������ߒ	f�����wv����|�^�)�8Yo���:o��d�κ��v�a�b�i���,Wo���/~`<Ɩ���C ��
FrmB�2_
?��#��nv��FM�k�����b�.i�%CT0�����L=���L�[PK�&'S��]l04��v��8/��z2�s��H4. zj�0������5k6�,"��6�q2!�P=<i
{>��2��K�ɑ�Ǫ��r������,���0���
O(��Q��9��N[]�l'����Pu��(�޽:��0�ZZ���W��b��#YF(%^���S��'����ܱ����̨�Ũ�)$y���S�8aH�3���9y$���j�>��������-�^��l��E�*D���a
σM���r����@��|uL�6��
#��I�s3������^%�ڸdiO�*�+���Л�P"c�Y��:!%S5�h��y���G��k�N5��&��f����i��1'z�`��
K��T�J�.W���p��ɿh�'�Q��]4k��f���Ua�KM�F+�Q���fYDW�*��c.�g�j��C�2,�\�z�����ǯ6��,�l��Ԟ1��N�j�ꓓ.�%��E�A��*�F��>*~����#��O���ݜ1�Pr��ϝ��*�Q2�H��x�!k"gw&7l�4�?̴�f�(l���iM9HS�������������K४��H$�u3J�%�W����Y-�Ǆ��O�G�R.�Gp���Z�V���S�M��Q�����8�gAM�#��
b�K~��Ϫ��@��6'�M��i�ٻ-eܳA�!��v�M)�����F�^?=/O��U�bгsY�]�y�=�"!8s��H �ԩ��J�¢���@��y�_b;���ͨ����mp	x}9�I�KO�KY���z�hᢪ�4�39/������U��aG�Nu.�տ����"��áJ�=�Pʹ��hO�Eد=��	
��L^���@;���k}��� �𷹻>5�~	��9Iz�s[J1Mn�N�b��M�I�ꅽu�c�ͦ�YH)�aTalb1Ůs�뺹Wc��5С��n����"��NL�EU� G:��y��=W��C7;���PS���).l��~��_�"���mx�扣ITyz��.m�4R���G^sa1��wm����:�p�M�>������NL�xѬ�|�S[XH��+&3G��k�g%1�n�m+�'���&;$���<�
>h?�R��Cm���r�U_&��o���D(h����ג�����(oT
���� ��v�B�_��(��q�.��0q1����L8fԍ���]=�ה�TWm����"�4��FJ�`Dx�7.�s���~Ú~��5BE�Ĭ�k���s+�n�^���G��q�+Cr�%;0�^H���ؠp�~]�R��ʗ�'����]���5@䃹V�Б����F��'O(z>�
(�z���) ��������P�j�=����OH�>h���al��1��vB�R�U�+~��4G��GUHK`ʹ|�/fe�m�_k[W(p�����̓L�)kwB+*s�WOd9�G�ؗ+_�g�1j�5a���`^B���^�rXko��@�T�e���83���.#����*�#4�;>&�^�Z
��O#���A�E|ns=z��"��������rGC�c���`����~{�����,���3�NY4�"�4$�A��l�.ʃfi���d~�i8~nD��F>�V[{F�LN��n�a �� ��L)":��R9�&Z��U'R