XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�I����QR
�0Anrl�%����_"�W|
��G�y�:&�D�o���H����!R4�I�f�yPnK���.�J0��Ε��!iXq
/5?��T�W���=m�:�/�C;�+z�x�g��y�4���3͟x^���/��s.Y�������%��J]B)��J�C�RpH�j���K���w^Ɂ����Zvb��`�֣α]�
�[�f��k[����o�( 8��������R(Xw����U������i����u���d~xL��h>�� ӄ���U?K�e�.�yz��+��d~�W��R�p5��C{���@ Ǔ��|�g?��P]O{7�4��J�,w����M����c��t�P��QH�&+<�c���ڋ�+��D�P�OG���>�]Xp��x�ЬĶNg��W�t�qɂ�TJ�m��$��?@�*�ɦ�������A��ϐE�7�t�uf>���w;�/f�xgJ&Y�v�_�'^�|�UXR>���2������I	�U��5�>W(L���QƟ��
�2�4��t��C4�Q�C��q\���A3q�ԩ�=vP��!�h�	�o^б&�`�Z}&�f#<u*"��>Q6*?{v?6�W��@�sqO�lڿX�e�'��Z��:�\ܚ'�ұ���k쇚˲r$�d��:�
�V���&�iY�$��r2��zܭ�����Tԩׅ��?�ˬ���vv�������cx�=k����vr�fǸ�=S���XlxVHYEB    b631    1a00�^�C�+�c��4��`E�:�Pu�t�Y��=���#C�1��TIa��I�8΁=�AWҩ��L�"K�#W���x ��N�N3hg���$�$bt�ݟߩқ����bU	X���{�5ˣ��'I��}��Ń2c�����R�+m�_G����F[����Qa�q�eP����O����^���y���G��\� �p���TѪϲ�^-#,���?�5�K�	��Kj��(jT�븅������>�mL�e���P�T�S���m��@F�i`-h�^J���Aԝ�4�Ɍ�#���gb�4ef�Oѽ`��g~����&Ҫ��R���Έ7-���Z�Q�	�x�������Ή3Q����$bʴ_�=�����=���v�S���V�SAg�oqe�$�R�k�R�̨��0h�-"��؜V�{��Y��AM�аvn,+=QNE:�A���^(�!V�tw�X2:kIGp����l�/�yY�\!<���=Y��`�"_���+$A�
�f!B�U�@$SN��)? a��2]��*i�r.=��텅����팠x_y喨e�%�z�om.w�ڨ�4�Ȱ�f���>� ��%��oˋ�]}���W�,C�޷)k�h3�D�gp&�x��x�*'�kWt�N�zJ�&B��}��mfر����ˋ�-�0ĕ�PybYDr5m�Q�zq��[�;���c�pUН��av��EYv�Ҙ���7�'G�OG��I�_S����3��cEF'��R{r���u w�9l���!
栤r�[�_�ͻ9!" �Q<�!*��<�nnMa7��q��<)S-?��^d��"����Y�����.:��8[.�4��Q�3�yGyg^	L��K�l?���R��3	�s�ޅ�ql�Y��r��s�е�_��~�9Q�HxKï���q|h���\���wn��'��S�Y_�����LFz�$��K@�kha�rt���~�����>�ի�N�-�B�p�L� ��ܛ�Z�
mܔ�S䎃}�k��N������[�D?�6���`�t�Fg�;S�E����.�8�j3j��	6��/��� eM6�Pn"#��E����,l���Q@y��^R��z��N'��g�k[�@W�l����|x�5�R?m�-�(�
�믇V߄� AN�a�dK�%�;t6l���O��Ͼ)�o�����ߺ��1Y�G�˗�$-�f��������p��B�lb�TL�Z���Z��X�vu!�����˗�	A�jc�EB0�����cc�|K5�3����7���/Z�L�'x�B:{�zIC]��8���Mf��6����F��E�^��1�nMsZ��T��Ӥ�3|C;vA�N"�X�&3��l�Y�>�4iH����
�P/Z�Vc_�a�Ϊ/�I��h�?��(}=�${gM�)���[Rn�<����,���]b�*��dy��}'��R�{-�J����w����w�6�W��S�q+n���5���Ma:��/�����E�M�܁���Q�h�vϫ�N@G�[�-��b:�	<�v����wD!���f�\ �u}�~����Q��d8n����k�Q� ���%�<?�'����3KK��s��̈1b$EЫ3�ڒ�C��M�P�omA��H'N�����3��/t��Z��?�/�o_����x���RDX�^	�OJ�Ϙ���؈��u_��'��-V)�	1�x��2~Le��Z�(f����a�O�\|5
�D�]�Ȍ��R�R�! q�ݷ�qqZN�FWM�7c�ʼ�9˗IƋ	�n�u��ۓ�=�&N�i��I�hDlя�s��+�6�H�c�Bчr�S�6,��mW��s��f��&��T@���D��wݰ����#�Z.�Cx�:t���	��(�	�"@���[���ÊGn���r�z�CD��}�lu��Z+��dQ��������h&O.���Z�_�?k!���b�[T��#�!�M娀D�p&π6�Y��͸PRD��L����<�OGf-<S�������k�1UG�'��5Th�Z֥�po
5�bx⮤��(pmD�a/�����SN�`3�/�t�zq滇�����^��	S]��@(V�>������DMù���B��0�����r����gY͍
_��*k�g�U��c��'�������,0�nQ��I�~��5�B��J���4��1'��u�cz������#��cJ�~p�kԫ���q�����zp�ؒрM��
�����D���"�����~�~ �j�qŖ��UJpaֵ����N,KN�q�=��'�`�����C�I�a?ńƢ_��B<���/>m.��d�M�Hp�JΆ��qi����
īK.Z"qh{"��_y��3�4�t� 'FRL�f�QȮ����Ԕ�2��T�v�Z=��O��v)P��8�2,��+ǿ��$X�Q�^���s��Y\[	
p"�E �Ձ���^��$sD�.�-���z0�Vο@����c�4��k�?�@�m�|b/��b�i��V�����z��Zi������8���d�SK��d�ĔL~�_7�h��JbNİ�� �#�ǹæ�jX�d`6�k�Z�h��+�ʒ9�R�|��5�_����9%����p� R�JZ\�1��f(�@_磩��9���'�>=_
���R@�U�F�[/����v--Ȓk���go7�:PV����D���9ރC�Y��)D����E���To�nĢ�^_w�mmo6�g�(��y���=|�������]�~�t��(
жLl\�C�Aps���Z}��h؃�P��1�r FZ���֝߹âK��-ݩ(�L�'TP�RE!�S쥒^��Z�.K�!�ӗ�O��J���6g_h	c�daZ��X=|(��]X�U� �圶G�s�_[\��.Z��"�Q^���Xa0PV�rs_��Tq&+���O[��)'b�"��#JM�D:�%L<�e��D*Gg� ��q�v�">bG����~�����w�Nd��@ s�kA���e�e�$�m���ߚ�_N�1��m߰V{�˴ݷ]�&(߅�e��Z7�+Gl���n��?�tCX���@ S�9���B�i��8��1�(��!��t�vF�"6����t�5I��!>�ƭB=EOmm-O�@|6&�+L C����vǔEuŔv��G��"|���� �ʹ� ��/$HC�Tz�ևH��M��xy�O&PU��	|�!�����?���J|�ݚd��\:|�t+�I۴��i��FCg��Hl12�)7.��d�� �7��1�@s睵�����Z{v��x�F�2a�h��.w�|�uJb�E9�����Y��?D��ibӖ��|�/<��!h\�t����$?]>'K�-�]�F>0K@��G�4���#��ɸCY�]kj:�RM��8M��AI�*�S�Z��A�p�GϜ��9W-�9���x*�&���,PK��b��Ax���}�d0`�-�6�"��(���.�xO�3��zqKN�e!�XTe� �R1f�K���Es�����zm��h���V1�=Ǩ����Ѫ,xXq�xb�X帹t�8! m1�kd]�ƍ��y�>VC/Q->���������.�qY�����
�����OPE4�6��T�Ӱ�2*�g�DS�-.��9��ufq�A���|ɤL�e8Nm�ڐ�];豲�D�	}�����3+���[�f����}�&|���R�{���Ѓ�I�j!����

wW���ht}�@2Ѣ�#C�}5����q�${���|�yo���Sݽ�Q4L��zG�y�gS��Q�Ġý|�m�N�~������9X�������Q�r����%���zY�h5�r2c��������{�����G�`͵�`�Ӵ����u��x�f�zX>�ڎ~N]T��}P�}4Ig�(k����P���q�M���7�C�#�
(��8�&f��l>r"ʺ�Š�=h�eHA�i���WϰVފ���
q�˕��$s����	��>EY�dܿ���.��_��x��ZA���l�ӣb_X�>��ТQ95���j9�u�?�fV/�����9��d������#���M��=ڛ��ޗmW=gr��	�1�9O�E��r�r����p�&4,v�b�1"�53�hɿ���G:W�vɤ|�$�|��$ѵ%�жM�:��&	�c;���������۾1߅�ǮA��y���㰦�oIXU6w]��O��0L'/l���#�$��k�*��N1�x\��`M�~�$e��/���A}%yB��C�PDi�BdqfG~V���?�.At�O>-fE'�:�UB^޻�3���[���zL��� [�0�Xl�#��ZE!#����3&"�qJDvyJ6��(EsE�{�V�wǢ��E�N�,������21�T�gL�BqA�,&����O�w��/�vWir�Eϔ]��4�1�t��E��Jf.B?t����
(��
�IK��H��1�Ć����&b��)"AĎ�ԁ(
%xO��p��0���r����o�y��Z�7>�����>�8��M�&�'�J��AMq��	�U���w�4����WhS,8џԣ�*;'��Y��*L�f���H��댨Y%i�'j/.eZ�\l��H^�|y�T���y��>����6}D���\�6[u!�"���q�aD9���j��X#�v9�R��)�]�r`�(�9jr�R����#��/_p��~�xi,�I�e]1��~�6W?x��K.S_�C��K����桼�_��i��GH�t��#U>�������ڍuKu�cnHs���P�M!V8�>henA/_���+8{�����S�A�I��n�F��e$�D��h/<�Ĭ���m�U��m,�oγ"EȘ{#]�n�����	�ᶼ�	 %�$HWț�ͶX�C������F��A4.8�cד�����[x��H����Mr���̫k���0պ?@���kM�z�����"�0�o�h���H;u���7^�`	�/�.3�G>.�:Z��P�\C=�"(V<?�K�R���Rd�ǶŒ����jI(˹��<:#w�lX/
6�/
{M�j�8B��&�����OՓ��G̰�1ǔs�wX�1iu�߫%���Q�,��a����S�ӽ��r���ػ�qcp'��y}�Ï2g~\Z�,�H�^>��4\��}Q����)U�}dp�H��pbEK�Y*����y5��(�|��3!հw��++�G�]Mڽ���]� �P�GJ"Ci֗	k���N�!Ì^�����ni�ֵ$��q��{���9��A:��o\�M��&�U:�iI+�{=%�1j&�_s(�oWZ�@��?��(�8s��s��,��Lѷ]�wd�����ʚ^C�Si5UY���'-F�?�0Lۄ6BR��}'��,~s1�,�]Ȫ��+���x�-DM�q�x�x}O��q"�8�tak��?�&�F���ag���H��߃�'<���_��7,`hg�rۄ��!I�͌�]��p���`�B����c��4R��<�s�S���	�be-�tR�':�l��|6V��?���'w;?%,&��{�����3a4�&�Z�p���@L���Y��N�8aJ������'�Π!�OQ�<۸��P�|��>��`�-M(d�vR4!�aƿ���c:��<�G1�����B���Eo"��:�ޕ]��L�,�]'�fGЌ�MAύ˶�2&MG�Q8ň!���^�#g�ނP=R�/�7�%����}Jl��u��;v�>��x���dNr��jd���<�%q��=y��R����.�LT.�"����ʥ��a��Hp���O]5vNN��ב�'��@��&W�7�`;/�m>̐��Ko��@�vH�B�'{���:��B"v��$G��:��kRa�*�G�ַ�wm���6rߜu]�!j\`�" �̞�V4�wN��ݳ�sGKg �����Ê�_+�7��`���mt3�őIB�:�Ds��0��f4x��1�f,�Ajↄ7���I�����s�VT6�f!wXL��U޶�,��9IY_�K� ���`�2��A��5��SLR#"��:iT�>Ա)f�,�����:���������e���E��Ho��g�I�r
"2չS���B�V�͂�G��]��t����@U�bX(%�.,F��պ4��\6P,@��"���������ΉEX1t����g��@��As_1֗x�`�l�H�|�ϲ���@ל�^��N�8�Hru�"i��7K��K}��QY��� <�O��t�wK�C(�z2L�^c-��+m�Yʟ܍A���f���K�ou,Zd%�Q��}��S_�*��o\�
C,/���g�3�V�O=?R���Fsb���&���}�u,G��c^Ǡ4��y)l����ա��J�:o��{$�������G9|~8�b�|-��M̈́�ǘ@��{q������W9d�ǡ
��$$�.z<�	��Z.�Xg��m�P��\��~��|�+G��^�-��&���vM�z�B��H���=�#�����c];~�j