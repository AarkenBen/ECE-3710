XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n�B�~fJ�K1��=Z OR�M���@f�lJ�5�X�L~�K ��Yw-"]#+�5-/]Y�p��.�}
g�ʓ	��aZ�恘���/Q+�!^�jT��nꈮń6������(	�D��I���}S�Xޤ�w��twvur:ݲ�'h�< ����ަ�sJ���5�ʍ' �Y0C�� ���|#3>��z�n&�p�j�uX���,��9D�WU�U�76����`-�2�~br�߾����y�-!��v�^�½�0������<E�"�+_�)ms�K�)�oOR��-�7fx��:����M�`қo�Z�|����/��^R�mGʥ f��m��"��@�'B�~�.�ǎ�ԓ����@���)���u>;��N�y'q��3� ���P�:qӝ��$�ӆ���6�,��q��˗�F���r�U
4̐2��s��v"1���*s�yS�����s�i�85�4��������S7��O���՞T���=1w��D��Ey��Y�f��dG�{גY��dj#Ǉ�]V�9#�j��,V�<�m�a��'���0M�+f�<�w'��_���.�vh��XZU)���O���Y=p�~(WJ��w���@�l"�BR�N:���7�B�^����8CG�N1p����Z��,��*c�JE2�[�VF�{��d#����Z�P��tI�+�<H�R�M�j6�0F��U���&��E��)
9⦐�.��B�|�ɣ�ٴ�H�XlxVHYEB    fa00    1ca0��R����5��g�)�3�y 9-[��a�asd�E��� ��pW=�i�D����<<����(~K���Nbk�@p(vbRS�ɻ�$�4i���|a�����Yܼ`��k�Ct�Z0b�BMR���D~ˍ�x����(�s}~��Sy.F>�$��<:�J�7L�΍�������'�X��8������*r�зV>wώNR7_��X��|����O���O�]4��K:e�1�JVa�1��xL5�=#\�ٜ�S�@y���.��/x}�V��)Rbl�%Ց@Wޱ:�~@U��<ֺ0~g����	'�;�7<|p\�Lד�"uu��#���@��z˿*�&�۠l�Qo$Q�H��4tOrI�\�vx��n3.l�w��y����bBk����g�:F%���@��{J�����q��#	������9�f��-�n�b�ȳ7MFWǵ�@���o�G��R���im�5��$�;;���$2��;��L�H�w�LE����BN����&a�>i�G�o��3��ƖO���#�kQ��$�,�Q��j�1ތY&����6S �������ܚ�}-F}0Lz�1��u�2���2)�m�*}�=�(OS�g}9�W�QZ�"�g��?���ޛ�﯄�ޕeb�TV#����0�TsY�V��0[�DAM��`����܍r ��p����}<	���'��y&�
�T��$�=�5�55�#1��B�V	0<� ���幜�ti�[�-\��?Yj�l��]DO{��?��Ĥg�,^Ќ��۞��ݝM¸>;	I0~N���,�?���]�_1��Nh�����~k��5xIP�I�y�'PZ�Q�z+�UYE:�H9q���7l�M��ޑ?ĄH�V3$٪?�n&� �|<��G�z~!xTk��75C�eR���v#Y�z��1R�(��m�˖o�.d �ڲp�3�{uɌE|�I�;��ߒ�}�7)J[s\�{U�[�YM�p��T�T#����&W#���V����y{G>*�#���Iza���xa^T#ߦ��
+}?e��,�+�����"yiND�:Eݛ�Jf����R�o)z	������m�x��k[�x�"_<�/�vA!%����Ҋ��������_q}ٖ`d6�y�C���j�v�,z�n������_�3�A��u!1���d5�J.��O`�$E�� ӽ\�p��_���͏
�u�:h�o'��K(���c��"��/��d*�șB �O�TLRR�qǞ�2
}@u������?X�`焌��9�w�x�!�S�7j�ֵ��k��c]0���U�Bȋ��h^�ѐ���jHĵk��ߟ;֋����\���w�{�-�d�;�]���:z��R���3y/oi����dR��U�S�~9򙏈ؘ˞����n�ڏ*;����H��q��]�D��`�WˤuS�I%�~^·$r[e��*a����X�^<��X�X2���6 �#�m����3*�W�^C�7�)�L�ר �'9	1���d���ՍH�M��il�I'�3"��2B1~�:cz������RM��i�����w!��ͺ��L,׽�����:����m�$��tB雞�Dw�}�]J��/)�KP�����ŷj�בwB�t?�T�X�&AMnx�oE$�@�׆��҅
�����T����O���u�������nqڦOv(U�.*�k���=	�虗�h���Nz%�}���ݟ��	��A.�Qg��z5�y�]4Zf8h�&�ݝN9R�{�v����黈�H��{���+#���N>�Ƴ����Vs[Ҁ�$!:�7;��zQ����Q��/�l�s��G��^t���p��A��0l�A���d_���ciT��Օ/�\�ڋw��-�ޓFy��J���J�(��� �t���i^�=�W6�B���6��T�^�2��F�L��w�0]�,���:��8�_$�s0ơ��W���bS~�1~im�H�(g%���ϻ�ͬ��b�;�F��8�6WJ�#Y���R'��1���l9�r�yGB�w r~ ��8�@>1Z_l�����!�t�����T��'��zgKu��X�4ߺWH�N�M��
I�U��v��i�q�����~$9f3�H]���׶��L�?�{��Pf2��5���B�lnD����?�֕(���N���4�B��T��x����x�Kj&�a��Ht7�_�p,�mc,l�喹Ȇ�n���+L6s��p�BFB0�J"}��e�7o=�,&}S8H�~TO�� ި��1.e0�I���V<e��	,H�3�d��wH?�V��:�u`�����zg�ݽ�R��	^X߿�j^�&���J|rj�'R�����&��"#��W��C1����
9����j��b8�7��R��ጦ������)��&��i�J"�{�ObU�G�xx�ޮ��H�w��i �gTm�I����[RZ�"�$f�l��P�!��6�ݞ��\y�y`�4k��=R�}j9Nq�e�mԝ$^��t)��sε,�z���ƱK��H��G^�7!�W����U��p�&����త"���.'�q'�u�
K��!��ŨO<�bL�F�1��H d�/�k�c��4�1	�q�p/��� $�i"	�rƏj�]b@FRL��G@��d�WFh�
�E��L���g@,�/��Lq-*Z��~}XiXn�(?O���%�%f�1���z�Z��}����N�]|��ӫ��t�ˍ/��J�4��$!�Ro���`��^�'�T~��i�0���#�֮~-bx
cyg�C�lR�G]�|u� #`&�@�
��t�,�l��:t1jE�+�:���(����z��]������S�N;G(����³�:�l��t,���O�$���	�xb=�%h�E��U���)��9��W��6���ӀP^�,�<g���7z���c[�]\{n�C=a��m���JڦQ��Қ�-q��2�T�Z�᛺]{_o��^��l)/j%5���,��Ԫn�0�j,��^����L@�Ӝ�B�D��&S�g6 P+ ^��[�wi�C�)�t�Jش��@;g��pe����x��g-�-�$s�V�z��`xm|QM<��p��.'O'H��BE8�֪�����A��t7y��6��Y�R	\��S���o����-�
,rs7��g?�ì�:Ѵ��lM��LW��X-�w�kn�:�B��5ߊ��&�W�Xm;b F��b[�CG�haU�UC��D���P��
'p�'Ƽ��A��jY.���Z����)���x$i�438���4FsT�n��̬b��!�2Ŭ�̐�9��]?�]N�E����d�;�Vq�m�H3��q��d�Һ����}��nI	��=4��^��_D����s�J�;�*S�b]G�?�2�l��L��~���T��j�{�*�W�kN>?� �\8�E�� �ݘ3�v|Aj��D0(����~�����@��K��ՁZ��-ׂe�H���ZZj�G|�2vrgC4�צ�����U�e���)hj���w��0�!��=)��	�!�5@�x~ʊ��W���u�O���:���>Ҫ)C��A �O\MK���D+��B��=�[(�ڛ<,��K����^T����w��Z���K�q�y� N�Ry������V�E���F�6�u!S�6�ъ��u�}ӽ��%�p�6�6��:�s`�&%AJP�_�x}H��L� �	lf P{�"z�gw=��C�֝�y������ӈ��ı��Z�*ñd��菾.^q6I@�?���8.�U�M�ƃ�RČ��������ǫ�'�/�x[���U�iR����ǧz����}����D�o��e(����AWn	�_C����D,������j�O!e'�#M.�_�3��Hu߆�ٛv�N�3���@ScP��G��dfɅ��Ut?�8�ĵ��=\���n��^��~�p� �ѩ��U���E)�UV����*�SǾ��٧�o�dњ��W��T\(�$䉸 Ǵ��=rA�跹Z*�
��5��\�R������CT,r�]�'�UrkZ̾���$�0<s^5�Z�T��/�[�R����k,����+����
�D�>Z[ʾ���B�D(UȊ�"��NA�O�|6ZxfN&�ʙ,��_��\'E�sS����9}����L���ˑ9©<�����A�\:d,��5�V�����=�g8/���I���/PT	��2 �(1�3%�;4)�)��,�.��lu{s5���}V�0��C:�R��*}��!��al8h��w��Ul��AkU�%�Bo���0*oQ!�L���2��m?��n��M�"��\�a�F�H�
y��cTx�Z�z�����7�t�qz���r�V������g�Vc�`�D�։���x�P]o��,�}�����5֐_#�a���O������c���pg[�;[Cd^��D쀗^_�0cx�d�?��Q�ȭ�r�΋��ꭚڀ}l�rf���ʒ��Eb*yhg�9ҽ�ǉqB�R�Z4��@Vm`[�H�C�886�����"^P��x!��^T}ގjȹ��Oԟ�Z=Q��a�¾�/��;h$S<�1ar`��9�i��I�ɺ��o}w�1��Gf�$���C�i�Ķ�$���x�!��(�:�)�6�aPo����Iu��i�F�B�/X����%�NB�m������9��֢7�P�K�z@6����iO�@�{a��� L���fY��3]����?	�7k���@H55�����.xk��t�M��w9� ��Kio�B��A��^�.d'cN, �nI����#�пs�$x|�.7�q&b�A�b�Zc�p�����#
)"����f��.]�����6��?-�{eܣ�����E"�\QR��9)���v�.����+�H������ϽH�����L�/�����Wqg1�;�U�ܫ�s�?k<(&W$@J%���z
F���[�_Z���G�P��75�܈Bm��9�ĩ"�je�pp��形K>y��e�W8���^^��;s+Oi����5m(F���FMoCW��á��s�ʎ��H�K��4��8Sa��9��8׏qͲ�ȏ�\"a7�H=��dy�"��s�X���� �w��\D_�v���o���V����JV����<���y��n3���&u�����: c�xC�9<�7i�xAo�~-�(�+f���~0XFP��Z�
��Hi�O˨��e�����M�!�4�Q��������-�w�ݑ�vqň��]�Y��s��J�}���w)�������4��Ќ?����w���_6k�R�Xz%כC���|\�|*e�7����q��(D �B���Dd�5=I��n��V�ƃ(������&a������X�ޮԻ(�vU��N�ω��[p�`��s�0���{�O�wA~���n�����eyh�h����_�� �gql���?Z1>�l�X�(�\��N�\$x�B��+Lh|�=1)C��E{d�G�G��B`q��)�A�κhuN�@�PC�$oTru��H�:E�8_�-�RM�� �����WGU�A��E�sb�>��֡bS������(l�4d0D��|�nd�BZV!�b������{c/�6}�!`:����"f�}Ox��Tm�(@OX�=�»�����:1@�|N46��ԁ+�簗R�Ϩ~͇�u<�X4��,s��^�~�tF���8���f�Ib�p?H�k��w�Hj?�IcO���~��-}x����������2�� �A�d~p���Y��jSHt��>��A�� (r"�'FvxM\����w�sA�:{A\�� #?=�7c|�E@���j�K���i|}�:О>�㠊�%��&�\��M���)��'^�s/ܧ��nt��I*��G��������bՌ�x6wU~�g��|�jb�0L��VL�s�u�l�*N�B2c{p��^��a¤���9c�=��(��E�`��&��WJh�?�w�`�9�~Db��A�&&~ܞ3�+��C�<Tᡒ���C�b�. �0��s����÷��:���&��@�������]�ߜ�5$< /T���F��mI�����a*�^Q�~(.��[��D��;#����* V�B\��� ���
�w��T��=��'C��AVD�1�ЄH�I�iHCG$̏*��DtMh7���כ	Y��������z���8�6��ƕ�K[�<iSdd�q�ŽSgw�t�IG*dK��
j�������ݎk3���5{g�?W���H;E�EF
��h����sT[����y��v#�\��I��SM߂'�9LZA�7:=�����#�#��K�*��
�]����Lx�x�Z���������vY#�^2L����s�����E�G�>Ц,'-���9w�yB�g�s�<i�M�R3��cAΟˤE��u[��9���@*ʜr˘EM"MK��d�d7��12䝚`#�����U��@ ͇��5lM~5�u(�L��2[ �+6u�^�{R
�4����7��1HĂ�{!v�t�ܪ1� �^�d�Ga�R�C�v��sV���!O<�����va��i!S(��X��9B���D��_��䌄Ս��O�N��@�`3,�wz���|d^�쬍²�|�H�,םoÆQ)����Ji�þD��eC6��b�54:� vzYS��G<� ��o\�GH�/���%�
�3Bh��P�cPD�����=[�|c�{���_H����d��{�C�����x��7N�28�pr���z�b�(-�l{�)ۍΤ*�l��}�f^�|��04��r&f�rq�G��WI��*F����qi��5���<H\9@��Ӣ�&�w�c:�D�MR�0&V�"Cu}|a���d������ Àh��{�M7I��� ��S�n�Y�@�j�.H������P���-�?��K�հtoA痰�^GD�����D�A��;��]����[����~���������z�z�&�� �e�����]����,���x�_�	T޴J=<�vb�
h�D�QlϢ���U�}\)B"��:'.<�����'�����k�otՁw׼X�]��������*���)-��iCd�TASXasO����O����=^y�	��W(�f0�־�̕�5\ ���e��hI;t�-i���N�D:�,Q������p��������XlxVHYEB    fa00     cf0{dWpɀ�V�@T���}]?
W㪎��_.Oc�ޜ�N �oe�5�ޯW�R�oY|�da �.������#
׉�W���3r.�@��6s%����HJVD �/Ѱ9�f5����+���X@�!N�W�Ki��]���	�}��Yd���I�塛��~��P�����>"�����I�I�
W����|J�N�wa�_���Ă�����N/�yD�<5ɭ��нXT��E�浅�� ���Í���)�l��R!�k��j�x�~�:���BP���(���;�%�=1���k��'��nNn����rN��g����H��MP~��� �-����HGG�"v+�Z¿�U����ֶpedI�*w0���O/:�E�=�'���|B��1�y�E��H5L�E�W�Z7�i_0���K����n���p��\[�啋���5�od����J��P���x��`6j���;�2�D�=�xBK�g\R�G�Zf!���sC ���oٺ#8h�oD����HZ��)��aa�dS���K�J���E�׹�[$�է��N���P��$��4��� �Y���gy���b#�%��M�*w�/�Y�~�Z�9~�6�;�m�m)tƩR�`�u�}��X]��7��	4ʍ�vg�����?�G-A�f�W*�<e��x:I�>ڵ�Aƺ4�M1��웈��x�K!3��C�gR��9���A�D?Nk��_kE�3�HGк����D�6��C5�Q������΀��$�Dc�/���̛~�-PĚ�0�F���V�@��]���~H��$&��ޕ����O&�wN, q9�y3%����ro���g���u֘AM��e�4At%I�ok���9{������s�M��V��]�Ҍ��n��V ���SH`���Z��M7�T�qD�c<P�!���+=�aG�Ȼ�x�
�V�~^��}h�詉	K�������-�y�aE�=�j�i�� D�$!�ѧgC5ɺ��ʒ��d�e}�Oʮ}��@B�)�A2m#�����п)���|n4mƛ��\ YP���N�)n��۰�	]�X��"+�&��ʨ3�� pQ���q�q�:���BGt��b���T�-�E �]��4�Y�&��arD���N�T��eJ��<���ƍޑt�R��It"z]����?��jl�R���ա�Rμ��%$����A+[}$�weջ��i�릮K��/cv�?<'�_����ǿ���쁯p��M;��a��x�� '�K�j��4lLܞ��5ȇ&pR]������uUB��K�O9^�ð�	�!*����
g#3R�X�{=��0�z�3�0�%�D�$��:��~Mсc4�M���Iy���S6��=&�3Q�
��͍`��-*_���=��-��mX�'1S]n��mؔ��Lt.�]NɇAf4bU�gǪi�����fOe
׶Zy�D��{GTS�G߬�D(� �_��?�[�E��ٖ4��A�Z����L�[
��.�D4	s)�.kZ��*��a�ߠ
Z�G������Cz.O�h5 �S�U@ �~��=�������/d��f/��h�|�w��1+�@*���ܖ�?��,��m��^_��M�1@�!pw�o�#�SS���'��S�"z'�W��j����i�ݡ��g���ާ���X�����)Wp�N9[���Ca1�N �GO�O?>P4d
���wni���[�oň��k/��~�c#R��;�����d�D�k�����9/%Q�ᓡ ��<�^,�&7:K"���ͥ&�v)$(�)�:r;�p�x�N�?U��30nc�:���*
,,�?�Jp���p�W���)�)W9�HV���u�._��
!]��u�:�
E��M�t�=5�љl�n�͝���<ڡ3��u��d�H�i��fҒ�W�3y��E
��tA�Q�Y��j!�I�u�ƓJ��q��R(OZ.��0����F����uK�X�e��?ʊ3�&�:�ע�(���6�ҍ��B���G�`�-tcx��&I$������k��i����#q��c'>�#I����N1)���u�ˑ�|����vU��#T���s���:7%�D˚��ɦ���X���Sb�i,�YAJ�S���'�?��a���c���Z��`�}�+@��2�bT't���z���n�8�L��o���cdۚ��Fպٽ�WSsuJ�´�h���뽪��q���|#2�A��'��c!�*K�)67�d{-�W�����<���R�T3����(�L�����;��p���^�@u��] �8�?i�������0�tC� .3����t�K����\�[%t�񍳌�{����1w�$5W�LP�����Ǯ✰����������BQZ��\�c�Ο�5uJ���2K��ȎA��B��W��c��6%�������O�;m_�XO�E�pd�I��(R;ۦ����f�Z�B�M�h�֨w������۩'�bJ�?�>�]�m��3�]���k�V4�v��U)��F�zV�q���H�Q ��m|:C������aW�I-vt���7�:i%f�x�.��\?oU�N(��u''/%���y_��!��;�y���H���y�+�C@Z�$pױbF��1!c�����K! �!���DX�i�r���H�#� V�w"�w����n�9Ihr����R�P+fy�٫���1r��@u�M#)�其v�x֡�6M�d*v*7�3�xs�H�?ο$&CQ��Ȏ�@L"To����7'����%p��2ۮ�O�-��8m-nѫ/^�Ҹ��־�>�Ǔ���]�>^��KnK��Ub`b�ݷ+�l�2� �ӓ?�?��{��/����ջt>�	���ȓC &��٠<�����"B�?���9�T�� M�~.O��c��ڎh�j&6E�4Th������2$��8�_��r���S���^i�Č��ڜ�dw��a��eR>�d}���Œȯ������&�e���/�b����{Ԭ�{���}���^�+wB�cst��D{�G���Y�|bWj��.qQ�dg��:?��kfvdC�=�"�)�U���w���d�c�^tjPh�'J���1�{ ��1	Vbo6ޫ\�s~���!�&7�+$��7���jpӞF;�8���6���E�c��Amth��-���V�.�#
ON���\�'�����߶39���+z{'�2��c�#1���TDy��L�J�{Mu��E)Pv7���8������v,x�sD��qC���ܗ��cXlxVHYEB    3981     4d0��
o��Ue[&<$�玥h��A�8��%�9�����ЖB1::�n�hX�����y��EBķ{{�����ī��X����禷'D�~�ы~tܿJ��k�1ζ�R�A&t�f�97 �+"�:%5W%���8���oF|d $�V���B-���Mǘ�]|�Jd��OW����≔�C#�.Pjo�(y�����&����fh���vD@��)\��9��0���6���":�v.G��T�+���M��%��e�$�����Y~��Q-���X�d���N���F YM~D��'	��;�I.ֹ��7�n>���
v�\����*�Z�ہ4��$oP~^�F���*	H.H�:z!��*�:<�s�����g��'�ιX�.�c�[��N��g���ϋ=1N�& r� �;�Z���5��D���z�����'���2�:��4Ŀ݊U6}R*nw��;
r�'�	�����%9�>�D杰��r�b���&3C��q�uH��?V�<��@�ܐ��C��x�eP��3e�v=yHau�H	m�R験^����nq�>
���˘�#�E7�[��~�q����)Ppp-(Ms�0M�x�:�p����2^���O�$3�6�����<�w���]�-z�C1����j�j���C�RZߤE��)���-���G���)�R
r�
��5����bk�4�Mi�xS�A	�����f�[!�S��0*�Ѫ뒎j��Tk���z����!'�+���@œ����O2�!W끵Ci�~c��+�0'���.̂=4��e樅DD�(g!��^&r �v������BY~{����*ք�>���BJ�� �=��	���������돼(���F��Msc{`G[u�wsݼޔ{�x#s^l�����V��ɀ��洸[³�8�C���WN'�W�i���{5Ơ��ǌ!��Ygת\I�r��x�4�TqM�:W��2Z�B+`�r��f�rA{b�'|�=�0�Q�K��&���߂jeu�m���W�%{9�'�ƙ����)(Q�,K�}�A�0�����Q/^&*��ءq�-�=
�RK�zQ�q�a�M:<W~�e��uА�[D��?"/&���אd ������!˅x��#�Oi�����<0����W+NMDSOX2鮒�ո���fu�l}cM�X��!r�+��N9������%�-����C^���j���Ƭ