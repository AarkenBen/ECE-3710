XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����IJm��}�pq#��،��ɱ�J1�Ί���i�߱���{$cK����3��!h"mK���SU���DRC�c�hJf�bY�0��e�Z2S.��t0!����S��>���c�M7Vk���٦�ݜ����Il�Ux*\;G	��/�� {1��/&�kv��|�	c�)GU���)����K,ٯc�P`5�wB1����O�-���GA�Z簾ġ�\ݧ�&����3�_>��4��d��������;���r��֑|l/���`�*�`��j{�Ί+���ٶ�&!�XY���T�Zě*���G�]���o����%����2�F�=N���:�صN�@T�i*�[ig�>l�'� ޯX��Zp=mY�����c��]X�|'eƴP�V�5����?ㄭv�=����>�9��0��eh鮙��;����ק��$��[-6ܘ�8)�jٴB�:<������#��Y�a>�}J�{�W�J7.s-�������:.�ъ�(�+�4��a{#Li��*�g#���[A1��?�������@Z������!󟋝�,�b1M�O��˻�)X루j��g�Ҫӛ�F-���e/�U�ɋ�+�3C�~EA��&�za�[q
�ba�0lE�s�C���0����(�V��8W��x;�	�� ��]B��{�~x�y�B$ޚ�ႉ��>����茢���ݴMP�I+/F|���-��g���-4T'{��q0 n�)���:���L���D-wSwG�&��XlxVHYEB    3042     c80L�Cfb���"�f3��}7��t���Hynl�x�[� ��qf����[��D��^�U���A���e��˯���,�7H�mB3=�x���K���B�@��W`�X�l�T2���F�~�|�="$����c O�Xl��s�Q�4�ёp2��t�'	����Ǩ���';'�l�319[ʆ��Y�t�>2^Dw��,��ϋ��xq镡�I�Bl���Iu`����	p�-�[�u�ڕ�y�om}�Fv��N�D͝��i���A���@q��X+�<O��R�L��Y8�L|S�^<6��1�R�<��6��n0���4F?��#�+�S
o�fN;�b�g��~.mw����Q�T�UW�yk�q������ķ��e�4d�r���Ϭ��w)	a�W�V b�&_���?����!�g��b�4aQ��QU�AN�s�I)�Ux������hn���Z-��o�
U =����v����@���͢2��{���s���Z�X�SO�����!����`,��Vs�����'��@�x���R�#�<�6ê�rb���Ӆ3n���]}�r�(>��}u�̂
P�U����Қ���B皩��o�փD���x)"O'�{��0ƛI~:Mj]�b����Qȣ&%�I�ę(���u{�MID�/f��;�mJ�WCx��x�6�T��$���7���@�-(�'�>:\�킴�1�!�\2h�þ�MR�棁>\�įd��cU� _�'n���ױ�-����:`�Ĉ�F��l��=P���k�
ę6��b�A�	أ����%� �����������ol}wT�q>1l֘OP@i	^�pp�Hn�-�~ |��0��O��6K�JBCgpN9Vi`˙LS���4�����.�OL���"��S�V��}�Q���B��o�[+������݃���>��.BV�:���	�_FM������|�h�o����X|:��������������zQ{![%.3����a��+����+A��]^�*�]�Az<�꛹ܴ�f���cT���E8;��άI�8�_��4|���Q��L@��M��%�+�tː����f�� ���M�3��B�����g
�b��>K�]�K�a����N�c���=cV���ʇ�r��e-Rh���/�!�E3�YM��p��y��z�|�8RQi��c�ł��zF���Ī��oH����� 3���HWA><��Y�埝�6se���Sh�H�+����3��ض��a6�'��]n4���H1ެ#�����H��w�)�3�m낛T�;�T�If:��Xx���]#hB�9y���&����N��q�
� =���X&-�l�w5jB~�0���EL��U_r���̴�f��)q#ͯ��<��6
�����yT�#�mݩi�4�IV��X�Q$Z*��>~�q�D5,�=��_�7�`�K�|,�����?
�Km,m��S�`�� ��oÕ����{�;)���8����4&��=�����G���m~]�*"��-eg~i��f��ʡ,�+��̒��<G�T�j�؄F\����������4����T�?�l}��!� DP��m,�@l��,�o����,����EbB������4���^� {���ǃL�dy��/*���ϧ�*g�����-N�/W��i�NA_��a����,��0���Ƚ�(��f���G�R䰔ؐ��������j7}E��5�Bt)G],�+ݟ|���̺����d7�����g�cU�$^�X��q����I�V�w�u��*�oOP����T�E� ��A�t��NOA81���2�)��?�l�;Cp�X��'�f���>��(���A���!����)��ƥ�i��g	�\�ôp�Y�Nd��!�\���j�^<(��n�E[y��v"�=J�Nxj3_(bˍ�#HA� [��Z#2l.���7�Oy�Yś�an.����_.#'���� ��- Vù��꛸������&ϲ���-��J=�z�p�S���؄�]O�ɞ_rWP.!�Ic�����i-�����U2|�S����֫oRV�Ü��<��5�RE��+�ЂBd�n�����b>�����F�\t��	�N=�N}V��_� !bع �L���L��g�G�u}�<���=Sq���n_��A��\��bl�K����>�e
�Y�%/�OQڵI@NO��&ƺu�5��v�;#!a �]�F���P�1�9Jp|�y��یq>�y��ʖf^�֮���,��Z�ɂI�𐞘Wz��v�=�n�X+����G�qo,- -ڛ3\��K��"1n��+N��!�Ε�Z(��*��>�]Y������B������IȐՉ������G��� �*�m�$��(r��奎���*^8�"BU��{�q�s�װ�:l&��e�	%��g�JV2a�c��g�USC媰��?��J�����!�hJ
~+%��bS�>On?�L�u��u��$����+qd�UREuP��wxӴ�WcO/��&w;�4{��ہ��+���n�N�����S�[i��� p.q��I��9eK.��Fjm��@���׽��3��0h�c��`���|]l��_���07t��&>�@�j��Y`��Q�o$xRFi�Q\f|u1%�T#"����Y��ꍢ^�۷s�n:�h����pcXN�$$���3��g�=}�z7�%YB����Ԕm����|v�#nz�I��	4[<�3�H8���3�SKu����)O�u�6���\퓍��>J���Ua�n�$�#��rȾ�M] ��5K�󰑊z�(�/wtt��Eq%q�l��-�yL� A�k��|�����ߣ��L��'FW�fy�+۰��o4�Ԩ�w)4U!����'�'(�"�7kLv���U���c3�B<���1fVSu(Z�"�'��:zX�Z��|��F��^/�Z�C̭*ހq�)�xE1Xb�Т&����!�p�~8Nk��(��4!t=.9��[C�8���s--��Ճ��s3%.�G�"���[F[������
rI+H����Z�Ld�ܰzn{�qylQ��#e:��r���2�csGț�r6��8�]!��ƚ�J�K