XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѱ=�|���;Sɀyܶ��~@[P��L��.F+�g�
ֺ8���a�Dw/�����fMM���mٴ�*uU7e�ɜ{1�vֿ��"��l��?~Zw��N^(v��Tt�T(�+�����u{Y�?�P8��,8�������Z��$?.������:C7o�4���.�^����{,?#9h)g��w��	��3��wN[ƈL�|�3�Êcp6���s�# �̓tc����T��Nf��L���*Rd���i�J;D;;�����QA��,~(��]��쓲HTX\r�.)����`P@��d�a��V#�\��~�I$���&�Z��?D>�"l9U<��Ί�+9�H����q@ْ8.�2���?�3t���S��F����&4oۧ��[��{c�/�>�Z���2&w�ze��|F�"�l���.Ŋ��ρɴ|�4�y�T����^Rw�q��x�MM�3���aMΙggG��~s�Sq>�%B���b��O�w?�;#a1�1������qJ�-���'pON�o��2ځ`�����f�ƴc ���A�O0��F�����i)ҧ�5./(d�M�)6BΟ���6���'$O�W��_5b���,yj��H���ʃ�>C?�=��9x+�W��iLp�R��	z�N��������1X<�(3�_���[�$�E�E��{$� �B��.�qz(����.����X�u��/�t�#"���k'�p� w@�4��:���,�X�"��}�fw%*XlxVHYEB    aa31    1e40!�<����g���F>mۅ����%~��W5���R%��9��g�Y�?(?�>뙡���i�85���Sq��b���9���Ji]��n$lO�-k����Gc��'��s�s�ڧˠh��p*ȶ��dc��3o�pC���u�mU���ɴ�A.�|����j�N�"lH+�$?̕W�5��x�X4��_fkl�֠YڴUe�1������{/(x��Arn���L0p���a�v�=����E»���0�ޓKL��˵4�B���P�w�_���GO�����7�-)�0O��]W����vs��<a�h�D�
�8��T����3Ga�eY��10-ق�C	pGó�遥 0	zo���� ���b�@f0�`5��ڳ��V��=�% *),bN�v�`�������4��pp"�q���W+J~��o=��,h���3���\;Hlր��C��M��Ub�W'��5��b�V�_�le�"��}��M�[z{!8=­]J�\�i���5�v?��+T��:U P��u�	�_h��Keux��g�K=��-B�\�brD�`-C���-m���!w8�k�{�P�S�EU�,1��ױ����`U�a�y*�u��1��n��FQ��8���\�+EC׷�E�#2O�Ǖ��x����p�ca��/	U�����3+'*��o [D0R��(lM�vx)*�e�ܧ�4C�y<	�׊���"�a�x'W8��:d�{>�HPP����z,+#Ba-t��C�y�AGI�/`�m�'q1���Ų�L�- ����<��H���6KZJ��*3�.�b�ZuO�X��pw+�����f��)ž�F�-���AM�X�Mw{Q{���}YL yV9ck}J�d����/��~����;�N+�s9�����w�
I���$p1?��ɸ���1[�����D&�6��&h�� 6��n��@�Y��Dڳ�,���h�v6�}��}fh�����+��@?r����\�����݁��#�Z��->��!~���g�J�ȱ׆�"f�B�(��;w����D�x�5�vI��V}G̦�9�_}s�	��+B���(�j[��$�ٶ+�K��>��h��Τh�k�J>ٰ=��~i�� tH[,��g��Z-Z�4�/����A� D��t/TȜvj��-�D/z|�KJ���	�I�����(�F����h���d��Ȧx{�x����s�[_[)�SI�#��f�C$u��fhc-,0]REHu>�K��Ѿ�6����������[�=�0�"���s]�̪Yj����1*Od.�i|{�J�c)rD���>и����ݮ�� �h�«��4���e���/���,�H�4�A�cP���`(�����E_�n��#tc�r���>��_�G��y����e�?2�^+����gV�jr�9�f_��iH7�*�3�A>�ZoLV�
��� ,bZ�#ASe�EЏ�ְ9$��9Ku9�L�l�z�`���%W�`�Յ�U��Y9,V�}��u
C��Y֋S?`7�63b�ԡq>��M���)_��y�C�$��Q�ٶ���8B	q�|�u�B0t-	�atA�Eg�3e�x�_����C x%�L؄�, ��o�M�*��EJ�2��c�^J�#��s�x8�O���.f��L�z��2�b�W�Q��C�U��&�����7��ƤJ��h��Q?�t��Vq�L��j��w_G*���͍�jV!��3�v�j^5�3�U��~*?����9��q  ���m�rRWy4�L�9_%8�!���+o�$��w]ºE�q]N�#m�u�q���� U��
Nbn���Jf�����+��:��@��N�V�A�k;,�iڠ_�h%�x�o1�)� pi�d����}�����<Ad~UKNc������)�cR��t�0�,�B����W�G���*�$��sy=�mcɆ���{`�[	E�@��{	P�!_&Sq��<NSOt�,RG�ݧ��v�&ޖA�G����VE5A��"w-��73�g3�6C�x��M���N2�ZJ���W����8U�9�o�'�l�k]8T�҃�PǑ��W�A�(s O�`��#{7�S<{���a:����?)���.^�P�d����W�>��]l1���bug'|�m��"-������!����0y�HW=�����wK��� �uD4��l����](�j7���Xh��ޖ7��Δ��:�/�$�B��V������Rؗ͠�q�� 1�g� M�B^{L����;N`�X�R #��Ը*�&�돸��8���] �(C,��U��+a �7�k�o([�ҿp�����9�Eu��0'�|��kb[��OS��,�)��5�B�hjl��p�.��%���97�Jn�,5��r�#�J���������ǔ��Z�����x�@}1j#J�mQ6�R��,5<j�Jtm�HcljVi���P� 60�V�:r&W��n*{�;~B�s���ϳ���d�27 �.x��cզj-͐�d��!<��v��5awZB ��\��%Wx%�`��u��o�������|(e�����W�YMVmG��7�CTmx$duo�V"��4�Oo(����z+l��'�ь���x�]��B�
��i�y$���I�<�q?�����3����' ��maR�> VL�o֤���dZ�QVH�	�Au�*����l�M�z-��oڝ�_7M��.�g��9��D��&��.Õ;Z�cg $�[���N�b��}�֙;���x�:$��Q+A4����Yk��-w����W���	�v��7�{^�@:����v	a�R9��q_�7�� ;��Hn�����@p����<�V��3��~�a�7}��n����<��*FP�t�@�҂�G
ݒ���;�m`L�qs_�B�2Qd�k�/�S!''x_���`��ܳ��Ӑ������h�^ �Q�tzz`���&��q���浲:=�T��0	"���~���E��~/���u��"9|�\*ʹ9�UAۏ�����nih�ￚ���|���/}�ҺZ�}��b�'HX�T�98� k�J|��T�����{	lAY�����X}Q$��|>l_��krX&J�4�Ĉ1�2Z�v�K����#�^S�O�H�/؟�d�r=�GxKsB� 7�	��oNJ>�G~B�J]�
c)��]wm�륏ￂ�;���T����:�)`�,����G���=��r���a���hQB����k#d �͍"���ݑ@57\�`�w������'���������)�^n���%-J����Ĵ��k����e���� ��x$CF�ormx�ԅ� v�6��'`��@�U�u�}�4	�pM].��E�[l�H.e��S��9B�y'͏e��?v5����9_�$����B{<���&��Α�t��lk	�LW�1���i�r*J3sD���k��3�&R�9x�C�a��L.KY����y�n�W��}h���`��4��d����Q獳+����g�6�.��G|���B,R���ΔkVJ���޶�D,�R|�yK��_���,���RS�1�{\X�t�E+h���O����X���;s�kv7bW�Y�o���r��k���M���T�au�Ox`�Yo�N���W�8����/����q[�c�g���o��E����g��?�z�vIz��P�\q��h-�Qb�_�'��Dԏ�"�g7Vo��]��ڨ���� ���y�`��u27������v��9v��J���z-�\�`�@�e��7��[Y��\���?��A�#����T����,�}���Hǲ�XtnƉ��	
�Ʒ��x����`0�K�&���?��H"������,��_\��vЄ�3��B�����Uh� 𺩙����;�m�,�G�BՅ���c���A��Ds��1E������ZgimGL��$�g:9��yF��A���?��r������G�G�0q|>�LZo�[�oA�G����2W�{)&|zhvvC�
�k%7��,����)���#��M*�~��C�*�i���z'���=�ARp��L��$*(&p�z�*��c��3-Ϡk�����:.�+�ð�7��nһ����b(�n��pl,�8z7�;����Cp�a9��/��u0���ΎU����N5KXĸ�ra�k����sC^��wtS7Zp4�}U�v�����J�Q�)Qr�],����0�Xn�9 �Y^��d2��?�g3ꔘ�Μ�B�(PC,1 �.���Mu�M�`������~��*j�ڇ�:�s��.�B,��7��c�=6�|(l7�[�brv�>�[�Rq���[g�����ҳ��
��jb�{�u�՞�y�u��Y�'I�c�=:M+1� Q'������6U��s0�%��,`/rCC"\-�G򳿵)�!<4'��*��.J���g�����q����!��`�"*U���Tv|�>{�9Z����b�oibb�o��~�4��閦��dQ���J�Nq��g��g��	� �y�oV��ϛ-f�����m�
���7���%ß��x�m�ݯl�w��I7��o+�]kг�$� G�eu�
��P�
��:��/�C��*��Z�2�Q=������%�~����B�4���9�e��c��6�[��m9Pp�pg��I����eQ4��G����A(�w�	��~b�{��;?�a�����5�
<yA�1�j��>>�nJ�	�q�6�NO�UΑ���Z̷�ͦ�.2�v�Y�s~����Ō�9�5�a��\�g�KjpC�:�K	v�eS��|�������v!�4�ǀ26z�E��>��!��6��dqG@ԭ��~y�<�Ş�����殻�A�QM��&��(�%��C�����L}��'D"�쒤��;��v
�������ܓU�f����΍�ɥ�t�lq�����Cp�#�k���8��Ry�����oM����ZAy%��7,�p�6��a����]]���H�]�������s�Պ��lOV��AO�n^-����톊�����{����!�vq>t�Э@�g��1ɧ��ڈ�~��I- PB7��vr��/�d'������?R�LC��~��o�G�Ɓ��Vr�t���D�mje87vu3��@��P�Cv=Q)�>B�i�O_A%;�f2:�i��,d���i�|!� �h�k��*�X�uZAp��D����PW�&\����Ls��lj�������Z���DgY�,�i\V�00��s�L�Ź8\�H}޻J��QA�vi�a?W�@�|I�T�3�g�Ũs>3&ã�9!_O�c�j���⢞�Yz� ��o�k����V� �-	���{�z���|ͮ�"��^��2��A����=CA�[���32�VHΊ
LwQ��cW�M�����
/�,%�#�+�&�K��cIiY�&F��S��)\�p`9*��:�-F�"�0T�|�������ۺ�x��'����֛�����Xl����xd�
Ϫ�"�ۮ0�WU^����ص�.Ho�^T�Ly�A�>���8z>� x�����t,�����C��Sf.?Ca`5��P����0&:���߹x���(=a�ݎ��<<v�,p�f3���}7���q>�X�����O���~���?�y�5���V�w���o1�n�1s��f�v�H��9҇LM�
�~F>�U�.v\�(��e���+#��~w��ep4d �uH'�0�8in2�w��^��0M7�v�εy��������H���ךƺ��ޕ�G6HL/\>#��٨�\���`$`s���}lZ�1���������u:���=�
�-�g|J��)�e��d��
���������Fp;�1�}��q�cCBy2�M�,�-QI�V^5��I���zV@G�����O�=U��3yQe�y�]Gx�T��y�-�^�,�%_"�qTlb��|r��)�=�珹��'̗D1j��)5&���}���:,�u]=���^�`3_��U�
B�jr��*z�1x� b\�OA\��RI�;�m�:�m�7��g*7ɛDkT ��'J����/�!��s�~�k���8f��S��B�x	"-hK�'��jt�(��x:�FW<�S�Hȸ��Fj�Z�I��}�s��,G#�Q�/7,s��`����.����r�C���
-ڪ�,���t"qc��¢s:Τ�*���B��4���|�gI�L��\�G�SLn��������>�6jY��
���(��� ����0�N�W�T��V#7\��lv�J��ML�����0�hm�0���;���U���#�슑5�)ڀ|��X�%462��P�f���.�Ǭ��E���I=����qn%ܷv'3l2W1�LS����Xn]b��g�O~^�@54�� ����AY�Î��;>�2A�=Lђ!8�r�l��YuK�W� ���Σ̢tCT>�#��5i��Ƞ��׭�d���/�������@�M\��9R��
��[�g�~��)ƘrE"m?��K�a���g�JB/�*�;2 ���{��P���*����3Ư�F[�3�G5�P<��
�9�����3RfM_�z����*����=�8(�`���Y��>߄�FC�W��d��0q����(������u���Y��T�p��J7�p&|―��l~+dҹ$CL<r}X�{��"#S���� ��<��Olbڷϝ�閗t��`I�W�Cѓ�~Y��}�6
��8KP֬�e,k>��-�Y�W���ߪ�c�n.*pS��[�N"��7�:m������ԫ=�+�+W��bZIoPA��P��~w�':8
C�"f���J=�u��m)�X�d�4���[����Q>K�ȝ�h�Hg�G��,}RkY "��
-"/ ��z��E���-%�l������+G��E+��?=#��h�V_�5M.���`�	ME�Z�*r ��X��I�8~�l�#7�+���ųO�
�@�,�,?-�ٗSo5�A,x��{mM�F�!E�!}��m�<�Q9*m�6!��j���Hj��hкcPj�m�^�[p�Nc�m��/%��y�G 3�(���� �+��]���a�EB=1�fB��0b�i�C�lF�$�'�Y9�QnrB����N�����A���A�v ���4���{t���'%���8��<�p���W�A�b�6D.�:?}zy;�,�o���nI��3�L���w"s�c6{!>���8��,���*�X���V]��}���i6��Ϧ�X9�5�8��xyr�T�2�!gr�e�G��̋2��4�F�o�pk�s�;.ia��K���� �L�.V� �kߎK<�f�.��3���W��%����-������1�	�~|��Z�V�,�xx}��=����,#k"6���Q)�\#���]��`N�p:����"AKz�\�a�g�K�K��-��B��0@��m��ê�S�,hA+rF�6�@�F�%�_�W�t� U/�4����u��R'���= P�|�e�R#��LA����`@�
����kt|�~#�I>ɀ�M�JI�H�)���N�.�<"*���6�P(���{��m<�57���Q�U��Kmn������ɀ���M9��>wȂ�^�]�ۭ5�