XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@����=��!�%�O�p�*H�M��kef���c�;���OEe�=�I�q�o����e k�I�4-�'5�ϯ����C,F4�c|�� }���Uc��n<�9�I��᝘B�ph�-�~eb��̢ʹ E���S�jo��
U�͊WJ��~����������,Fn�57h���	��O����^�����E�&2;G�l��sԻ�L��b��h����;GƇN<ҟCa�3�@��D2y��v�t@�2@���c���:]�0�ɦ�ⶦL��j��� �̡�����n]�#���$8��O��J����������A��e%�k�m����)����~	�$G�)}D���q�A!M���0�����@~�:[���<�G)���H�(�
Z2����V�R������o{
��g#�<�?M�;5̊I�����$�
�޽���b�F�֌j�����c}�%�9Ԇ��:a�Z*�@��=g�&�Z�/�?��nWsd�WJ�+R��d@0e��_`����i�h�ˮN]~*~���������H�����t�ʁU�bģ���1�$�ͥ&�����Y4F�M�/sf�Q��R ��U�0(/��y�Z�w��U:7���m��٦{�pDL+҈.i��m�6��f՛N�e�|��-�����+��X��j�1��!X{:�������΄FFڮP���)a1BC�C����gÎ�X�ؗ?�A����^C8�6��J(ke2fT��&�~W��_�XlxVHYEB    fa00    2560:ƪ�J�(N���~��~φ���O��jªEf�~����|>c׫"Bճ��+T)�9L��"l*N�+��A�}�<�ġ7-��&fImsM�Ug���itj�����5\ǹ�RL��j%:��d��l��س]3�̱XDG\�1�*��u����\�����R��髖�m-GU�/P���W��qD�z�IG�����3�+̓��zF
8b_:�k�-G����� .�=,7��)a8'�H4G}pJ\�T/�ޞ��r?��h�D��=U<�ہ��A�mO����[�z`#"�m3e��>46d2��	�9sH%s+铍o�w5�m��d#�H��a�3�C�'^�@.�Rlpk�ȃ l�T2x�3X��g� o�� ��C�)I4[4�Fۃ�8�`r��]�߶�Cj5lT\�_aU����x���6M�����zt.����d�r��b���&C�r�� AƘ�`4���ߔ�1 2 �3N�e4�E(&8��L��NE��p���Xrb$ڋ ��������K"�e:C�'t'�]�3q�`��7$���a���O�~|�������]��0P��=-)�U%�	SF�	CE >M�9,��� �9�D�Zf9+��,o��|(�c��m�u�ڳxTNG��h�����X�����|����}��Z	�B/XKȒ� ,��U@؇�^�Vo��(y���&��͚`�\Z��c)�vG�W�9
�e����P���Fi����P�����UX��<��Vp�XC��r_�������k{cy´�쒬��p�E{8)��ߟ��E�M|�̇䏫�������5'0�����.[%�h�n����i��]7f)�k�[��Ɵ�E��4|���@G�$�򩑈>��Z.�?�+heg��|S)�#)�����<� pw�#c��-m&�{ߓ��aSZ,��HNħ2�����bE�!gò��VD�?
���Η��[Kq�3 (IetǪ�������ϔ���lX7ãC�@����|���`5�i�}W��,�c�(N�eE���c�Ő�@�a��xܲ!!s���"��rD~�H�1�~��%R{$C�Њ��� 3��@��'���@0��ܭB�iI_|з��|�L9���8"j���|�౾h|�S�����*�fό�&����J�{	,I�wQ��3��-�mw8�{�7Zm�H����*�&ٍG:�zݶ�[m]�*�c�{��C�|��`sL9�)��7TFE���>�P*/p��S��lΡ���[K(��#rB���3�������t��|Ys��)�߈J���Q�Ò铂o�Fx�ؿ�����B���W8m!���%�v�Ď�"͎Ur����tF��sŽ�D<C�LpK�<w{7Wkm��������ִg��H@z���}�|I�1��F90�3�|���|x��T
/��ʄ���>Qe�#aC&�J�a@�����/q�-ڪwSo��5+5��(�bN��"��Rs����Rdp�
��ƬMi�Pe:��X�y��Z�O��Tw�h��}g�F݃y$��T_ڃ�F�*��Lj��b�ʿ��
����@�FS!wcQ�k�g����"FC�jyӝߜ��%1��K�!Xm|CF���g���A�A�&mX�0PeH#��X�N*班14�J�k���T�ɐoa�VT+F-1���ѱ�Ή�M��	F���wȲ��E����UP�	^|���<���6%�3����Y4n��QP�_g�3����k��c��l����B'�?��w8�
T\P���t����[l�L��`��]��&�m�
�(��f;�)5zr�A ��>��f>)����͙R?D�~<^qM�C�:޲���4ۮ� ��e���ڧ ��ک���1vx�\�g�@��B���4��hq�\��8�����F�CY�N�e6qJ������vؖ� �0Jх[g?�Ů�BP>����"��3�p5bFn >�HJv��٫2�hߢ�&#�y�b'x�V
QE�z�8�ᐑ��o���aZ ���8�@�F�nO����A�xZ��OA�H����`�9�1�9���5��N�������" ��L'%��(�m�� �vƮ��c�}e�4��t���y��c�q�j�(���vi�vy��5[����7����\e��;�z�������L}f�����s��cX��k8xk����q����^����l�� Θ� ݽ��P\�����Cy)q%����
���>y>�̐�p3RI��n�7*��E�N��P���ߓ7\#�ǿ=��cӠ�Q�o�\����R@A�S��6��0]cа����8���4�ޯ����W�'�
���\i��J��nRn\����T�M���վ�kc��z�'ɴm��V1�@+��G1��B��ۄN�\B���6J����Ya�^-��hu�r
�����Ё}�y�cn\���!Οp�\�v��f��fl��8����v=N֑���6�h&5_�m�'���H�^W0{�=m��k���7�6t��X`$�v8��rrS�9��V8lp�D��QoH��)9^���.�,{V����4��U5~��������/	���4&ύ&�'����
�\LtH�a����z�; G�7�EG ����9DJO��?ֿ����L&����A?�������D��>F%O�LNlH_>����u��/$eC��������X��7zd�R�1��E$���v�(8�f���Lgܖ�湬���C W46�z����-@��K����W�t�O�^�i�-�d�^��?��M��L��B�B�7�VҔ䜲�F{��.�9�rJzML���� u��_���T�/B�5�m�Ŀq�ɮ��ӘT�TK�Ju�x;�tLX���[�>��Hm'ha�݄25%'����*g�)^],��r��u
�m�^{l�����qK㯐� (T/���]����g%��o݉͑s%��yi��]Ut�gs\� r��_Ev/A-�B�r�"�"[.�>��2	a���_��~���m���L��R8n�-�ń�"x�_<s��`�ix���t?д���C��پ��W+��	�\������4V �(E�[�����~L�����'b��1@�m�..c����\�Ld�8I�.��<m�vV��
m����,4:Z�l1�TM5��5е���DZG�����ĵ�]��A����K΢E�@�ԋ
�xVm�#�x؀�g��$�tM���J��މ 
�E�6��k
)�x���D%c�� b�Fz^ ���T[L�ǡ~�ِ��V4��4��N�z}��I;A�t��&`;� �d۰l����c���v�v�,�R~�3C�k�s���~�N��l��?W\6�RU�E;+��kj+���D/@���e!l_ N�?�]@]�����I+����>�Q�{F�	��{P�=�iqr�Ʈ��`��m�{��y��D�Ha�E*���jnP�޹�X�s��Y��Z['��]�BfJ���&���2FRp����y�g}���u6n���w���+�m�FH�3\�#��D1�"���i͋�0������d{z��O�
W��A}���
H���396 d-X*gG��D�	��O�c���GŚ�o&%�@��%L#M�{�1�Ҏ��+x-�]��O��@w�8��'`:�\-��{�m�H�¹��x��MJ ��'���a����kʆ���G ��ϲ1j��y
���&əۥ�|L��c�Q���t�*�����783r��e��.���#�h:��� ��(v �W��"(��-s1:gn�����>1�[�����hp����l_��zԋ=�E�a���n�!�ٵ�^rG��Gq;$@�U"�N`i�%	�!V�Z:�� �?���˪��-p����F=��A�����׫ν�o���?�����B�1�)�:=ל��&yߝ��2'et�(ږ�?A��{r��0'���bj_uԩ��9�]p�;��1 ��i�^B}����9��+W:Y?���2,QF��U��b�7�\>
���k�j(F��י˖��,*��vp�R��c�f5[����1�PXleT�B]�?.[�����1~nDI8@��� �~q�P�+M�lVi|�e	B=uu`��Q?�l9��Z*�����VOs��+��𿫜/^��X�&O:a�j�1Ef����}��CWͪ�=�����(J�S�Ky3��U��MQ�F�0�X!�Y�렖J��kK�$��t�3�?�N�@.G	=�-�(�{�+�s���V�|����P풆$��9�p~�~�U�gR������T'�
2@ȃi�8��r��P���D��:�{o�Z:�g z��'ݿ��ٟL�7e��'�]"���}���7*ҕ���_�#��|Aԕ�w����Lj5XBe�
G��=�{[Wd((:4�A:=}yu�o�A���E5$���#�M *����\���=�L���n�a�����r���7l������,���
��s����x�SÃB:��|gK ;�$JO��m�R�(��1u��NEZʲ����l��}#z}u�nE�6�k�]b�4�+����I�����ͬ.HKgt�l���V���:�,���$�|�nm�>M[���$4SD3�|���t�v���F���{0s䣛��[����l���4��'t��2�}�{O���7ae���M��|�����S`u�_ET��ڗ�J�6������Z�"@T�n�Eu0	��V��J��D�TU�����d���]� Pvŏ�6�����
>����I	�lL=�~5Uy}9���搨����O[C����,�-�|gT����i{	�)�FJl0����	r�w�u �m��SA�����ߢm�f���I��z�pyW�,�%S��#������V]�C=n���p`㯹_�3� �뿐dȅŁ��	h�_q���4t(A�y"3�j�GfW��������cG��h���n}�xA5���G��I�v�� 4p�г��Y�V�vܴ�" �w)"��B^Q`��`o�ؑZ�!����ɭ��N���'Y<����>Xj=_~	���w������? ۟��P�m�u�����!���<%�� �KB���ab|�����@b���Hi����S��3���o�0���h�.�Ay��Oմ�-�GgpM�}�r	�Dҹ����N��c&K?����([��h�v���)�:�8z:B��V6�{�a��ys$UE��Ȑ��9-@���v��V��|�L6�Vz�ח���j�	�����j/[����r$�b���x��|xV>+|1�%V(Ě&��[��Pa�&NGp�u��/����X�麑Wv79������S@L��/t����Wb����nx�o�B_�O�@	�U����g�� =Ԙ��s�nxC��]3'i?;V�7�dΏKRHa����0Kg��\2cK���Mk���'&��X�8���|�Pq	����|��r-��[Xk��46�~e�Y��E����;h��<#���gJ;���7$��K`�i1�yb�HoR����HI�IǤaZ�ep"Ѱ|�	u�S�p$5 �F�\�슚#�E�V�aߒ��Q+v��H.�s������_SQ�[�b��{óp�6��`���M�Jrj���S�Y�%rA�i�z�cJ�+m	92��]���< ��2�=��O� 8�'8� �6��}��V�q*�?�{L˙q����c���i���
�$�T�Z��qT%+YU|6�zxD��`e����(��7h��/ c��G-N�j����Sv�'kq�%i o��?�W��h��_'cC�.rKPl��0t�
�>��6�YOqb�?4�j����=�%0���>I,�Z��O�C�}�[r�X�z�X���16��������(W� �?�	����GL!��b75L��ByQ�2��v�.��۱�P�s_e]����8�;\��p�2|���j#9Ք�x �=#6��5f}����2I�ex�F��`�KV�t)0!cIF�NY����]�v0�6=ܦg�Cu��Xn(؂�
�:,s}�A6w皰����E�O��(��Rَ��=^��b�Ӄ�RG��02��|^y�g&�ፂc��/��׺'��D�Zp`��9E�>0%T&I����ܪ�CI+`��ҡ=�l��������O8}bN��t��I���5 x�G-Uw��Q2�d1�w�;��TwTն�H`R�iǢ��N��!H$k"Qq���OQ�Ч��1� ����Y�Nj�i�i�o�J��YU8���K�W<�^�u�2m^�0�kFE���(�:��eD������L�� �p���e䘳&RK�H!FU�o����A���=���V���>{��F�#̢Y`�̿��[	����6�� �Ԕ�*�����t�}f��C�w�9	���|�>^�_�!"|�k����QE�S^z6j`��2�>7�R���8X��в��r������
��A����\E��(}2�_����`fO%m��f�԰�������.X���th^���Tx+P<�Uf�ޤհrx#�p?�Pz���~Tl��y=�L����Kx:!6�6�n�*^�"0Y����6Ϲ��n�.ie_�TM��ޝ���K��L�7��qI��क़�T)}�Ȏ����Y�adfM��r��H�O�:�*Y)k���_5���X�DxR{���N���mp��^G"�I�neX�;T���d|܅J��4Q�L�l#�R���V�=��6�+p�Lk�^�gܸ�1�zߑCM�k������	�9�<��D�gz�,a���n�*���@q�����?��]z����Qd�&�g=��p��h��io6��S��3�&�����0\�DN���%�t��	W��^L8[=Igh�ll�YUS(������(�=�s�4ˏ�#V?��}�O�N�م����`��q�"�r��<��W��;j}�5�f�V��GA�6���">��
3p�"�Z��_�6��H3�$��|�0����F�<7����Ixø[�T�S:��G�SA�x�Jv�~�I`1Y�,��o'i�^@�kћ�Ͻ��}�?ۄ&>m�$���� ً8��ӷ�*����	ĳbډ}�ng��1� �v�!u�R���M��%��_vu��\#J�C��!�S�+�m��v�����;�+�-K!�.��?M��w�������\�X�v����_Ż��x���c�A��e�h�َ,����MK�6��>��GpP���V�C���L�e���z���2�:]�c���\��D�8�K�����l�"R]xj�=�]��虡 8Y��%q{@K3����?���c�^B�*?��G|Ӑ��ɵӂ�Nx�e'�д�ɣ5^�یaE�[�U)4㶎:G�_;��#5�'k�ǈ�+�Y]|�{������S+�p�&������{@j����_֙�責Ka��?7�<�?�/��Lx�C:T�P����������v���A��5�PH/E6DE+��N���G̪Q���M���4��R�H��WʘC|��gcM�r).�j����_7l�M����aCb?_K >�sX
�{7��S2���_Q	�f�gbW���6Hi��`t��Й�a����|;R���[G�z�,X7�$�U5r*�ܷ�V�	q��̆+�����j��s�=�d�E�C]u����i�Z�;�����Wc}�Ծ#�{ @�p�/��0�$��"��m�P�l�� �]8ԠLz�2�/�R'*�z��ѧ��u�Č�.��P�1�z3������R�{\�i(F{Y�-R��v���P�g�<�AG���$o�KD*��a��\nwBF�LGA�FJ�;���q͏D��V.����h�3��y��Ѕ9(ڹ���ͩkt�3�{jTI^����/lՈy��1D����c��1]�(� Ɠ2��Pq�l,��(n��k�V�z�Z�I�B�"���9���H�oťF�l7�����ի��z�����u�E�-B>�`.����8��g��j�'3��U�s�$-���Ζ���mE��ZQ V�
�DbEGP�o$\=���`D=�}��Q��fs:��RL�sފ�h�������0c�;��Sw��ݦ썇�0PCi��6�{a���Y|��%�=a���ZҡsV�q�����-�N���ڍO���/������#� lk�4y�����c�jIY�!�
yQf!1�U�DC-�;�S�2�k,�w�{ݳt38���.W�1PA`9
�ᣎN�t��n�Mr�tg&�p\�r`����l�3c�(:���n�M�:��R5�pD�<un��#�OQ"���qC��W	�.�)��#��Oaz�������ܽ,̓bk,l�a���G����%���`.2�m����E�c4��3������n��*2�MMB�Ti�S�A
o�O��L�t�&:�P&��<@�1������N1�2�JC\��ˏ9�cs�aڳq����<�w� ks�o�K8��~��T����I!��\��F�A�թ��
��.�.�tS��Q����I8�AO������_���d+L�A}�z�<z�\-�u��!!i=B�MIá!��W����5G�L�!:�Hœ9]��	�\=a?x��;���ԃt5�b��]lEC�u+���r�7�:�t��e(��N]Ao�'� JG&�԰�]8�]��U�05����O1�����K�|�h/�3��Q��S��n�p�~���Q����FW����az8X�I��ie_��gCp����i�;4��o�ŭ����}�9�
�۞�S����('j�pyy�N�F��Wx2RG���ÍFRltFg��B�x[8X��x��T��̼|(=�w�����:�o��H�����7��w>D�4�Z'G�΅�r�<�0?�#�1���GDn�r�	����J.q��=n�a�e��Qe��̴�Ba�I\YI�
��b[���`�gz���B�k�|��;��Kk ��JY���)�\t��K���X7�\�M_E?ң(8����)}����;{u/�k(Ͽ'�y�2�Q}�CU����,�
��=���S njL�J�s����Ɓ��2��H�#�����V�?����@�S=��@���rCn�w���iȄ�jm�^���&�8�!�v�mq�;�~,�l���QZ,��ڽ�N����`���r6B� ɡ�*u<�P��R��� �w'�����r{�
�v���&�o�6l����l/���O�W���7�=�!�������x��߹�_��N�-��o����0�7��������G��(�P�&�{���XlxVHYEB    fa00    14b0�iҧ�c)!��EޓD� �ءW6��vv��F�Kv5⽌C��u���B:��H�|����]r��Ȼ/�������$�tץ�{ypa9��xu4ʡ��kꄃ�c�o��J���~Q��ϣ@]T���%�%M�9���Xˋ(�u�c��0�&Q��� Y:���t^��N34�/l��O�q?�&�Z��-\��*%}���?�����_���E��\���jj%ӝm�G�t{�@���: v�D�{۝�=BGΡ��絘y�R\@�4����>S��Ey����;��W����������Ĳ��px8�fٚ y3���1���mM!?��݄�|G�O5�݋je*rz��(�.�ʱ�=_-�[�Y(0 ��^���[Jڊ���p�#�l��.��q��X�ț��<���v���G;�!���DU\�5R����7�|���ߩ}8ힲz�k����<��츳�V�T'N��xy����/<�B�w2Pz��s@�t��-/��X�T��^�7D\�0GW%M�5 ��U;��F}���yn^�|NFW��h����d�+�I
O�)Z��Td^���0�U:�<F�	��2��p�n?)�r��g�>Os9�K3���7���z���&�tZ�4���UaHH���cȳ���(�i��,Jq� e���������Y��״�V�m�n��l)��?��\Y2b�>Yhr����ߓX�LE���fR�"�����Z�Dm���Ģ
�`�
�vq#��u�<�����s(���F-�.���p�1��b�F�I�ٱp��⓭A���JT���D�f�__����؊���W.��0��Cþ���Bջ��&�Z����Þ���s�鹬���ʔ5�q�j*��Fs.i�}DDb,��r 0-�v�w�-��沖�C�I�wv��=	 e�� �F�X�ْ8�p��RۮM�OB�]�����`.. �d�-��+v/�jٮhoGU�Fҵ��C���s�w��*qas��e�e��mw�M��S7�^ֻp���ݺ=tm������DK��Ip���o��+
�b��`����A�q�%���y���,?�a�h��
�o2e�>��]�Z�%�WO��eFf?������ׁo�V���sC�oIL%�*eD�)p�;�<�T��9�[y�of�L*�����N�WЉc���E��F3�0xV�5�B��/E��=��(9��p �t��7��>�0�3��<��)�����p��XԥO�P��G����u�9O����{1/�ulK��4�p���&���7�_iWv>��
�|��������� ���粢��'���s�%G0��ls*l��ZJ���9{��}R�F�Ld6����n���5�ڙkP��6T�9� ���,'�l�9a�+�@7�n)�p~,.�~A��vͥ,TpN6q�2�7�AF~Ͷ>1J�P4ԡ��Y-�%j,tӨ���^�@2k�|q���G̸~��cOɁ��"�D�v�����H�z?g̰�����c��i;X�a�?i]_`�~~N2���:��8���֎��2�G�|��s��:�mX3���%��X�KYǒ���6������4�i��j�ْ_	���'{��=#��i7|X��Y㨸7Ju��S��d;�q�汮���~C����ER;G8s]��Tg+tM�b�L��;Y%I�� $
�pDVC�D:�+�ZF�0�4�@���NEv���ʃ�MEu����'�m�衆�wN�5��X�?��4�z���ͣ�F�*�.�9��gN6��/�u�b� X]yx���F��~ֵυB�m���7�
�6�~�r(� ��ٿ�6��-�p$"�O�06IQ�f����N�dC^�ԋ����h���<Z��>g�ѻ�i9�Yv�t|JM��0��6mN�$��4S������;��oq�7���wT���H��ԇ"���ܩ�c�+���Ru4A�Y �J%��W�y񴋝k�R]��fz�ʊ`�Ś�z�s� ��k5__Y$�6��9�F�j�b�t�@�jq�yWr;��P����3�R�K���/X|�ζ��U���NAc�����T>��I�5�3��YL�I�H�_j���e�Ru	f25�G���y�'G�R�A����q����v���ρ3�� ���M�6J'�����
<�Ѱ]��6��#2�m�(ہ�4��Da�F�&T�xۊHc����&kKv�b�&��D�#�*T�a���(Y�A�5�=�
Rrt�=7���#FG(g�������8�B�#wɝھx�l�:��A<]��/А<���-�?�:��h�_[>G��F�������uY�[�������6fMw�����+I���\���{)\z�������OkB���@(#?��}��󁓞a;ڱ/��/���cԂp��3r�#gjM(��v�5ֈvV�H���]Ͻv��\Wm�J�Ek�D�����B��;^�}�P:ro\$�IYOj���@ς�r۞&+�Gɥ	�f�;�?TӀ{��=�6f@����{�iVt0$�Ov���������{���iG�t�!�$]�0�k�=!v��
o6<���y�x�<������_��QR$g�C�3�����3n���邿Y:���V"ӡH:��X�u��i�1"Z�����v�
��풀~p��0���wߧ�{��|�����G��[�|��9���7޼��c*#p2z�0���{dn��qp6�";���a���j�B�e����FJpk��F������	�z��d�����u�r��ߞ_�T��H���� ST�6��3�uۚ��n���^�k�������Օ?��%*\�i�r񴩜�FbԮ��q�\�|�"u�#<l��/��H2PbY��x
�]�L����/�>�OEA@:-n!N��;0�1��K��Ɏ ���c�GF67�D��h�a����RܰF�^����A������O�Րź�Y�&笽�;�s%o)�_��x(}PAϹ��P0Zћj��Β�]ڤ�2���4��F�<�����3����:�~8�Vm�p4�:�!�j{!#9�3��l�:.���&���8�5�~�1N��������4�Tя:d��jYO�w�h�T�h���d����K�b"��J���i�6��g���N������ſ��iͩ��/��x@�����n��w�����~/#�l/�R��EL�'@�x�8�赱bF�0O%w�l�Дs����
rH_���U���r=���h��Hy��zT����/g�L���SG*S�ZK��}j)�B��\kx�b��W�ǹ�F٫�ڟz�	����3�G7bv��]}8�]�;@����O����!R#�t_Cb��k�[���qY�/J�/k�܊L��c���S���uJ��O64�3Fv��P�Iݥ��=w�� ��Ӛ�;�I,���	`�C0-�m$������m���ƶa5�j�2-��pb��c��GT��'9��*��6x=̗�ȶ��p�]O�i�o؀4�Q�w���bd��6�{�����$�'�����K�ԊR6,�ǫԒ/g��4�}`�T������P��M'a����>i�,q�I>�3���'���.�<�$��A��)�nu��omk�Ma����Ϊ����HW�!8����C�u%�����TX5��W=�?�Z�A����8p?@�I�����߸nڑ�B?H��!�
6i��s[Z�-����g��q�i��8��<-@�s���@���A���p����k�TƜ�* �}HDa÷'�b�v�����bx��twC$dM"dЮ��G4�w�\"ߕ�ڌ�R�ٰK����Z�kS�LYC���g��e�Zǩ4sv�&�fB���]�$`��������ؽ'�-�%�	8�@눈��/i����^ƣ�G��ki`�.ph�'�i�\�,l�F�z�Pu�i��BB;Z�ܧ�]�-gt�T��h���'���q�0 �f�$r���̥M٫�|�'���Yb(l>���I4\)Ɇ%��w��U�q<t�%��_70�'׈U֓.2��lB�JA[0,C��z�;�o���5�G{lb�:"5Ghh)7zo����t\��2:8������!u�-7��d��\�#1z*�K�̞	�uD�!��_{@��7q|�؇uI���j9��Z`;���gW�����/-[�����P=��,�x�NncY��=�qM�ނ%��Zɀ���P ˱��@���5ax6)��QY�l�&��J���5���%�6��Q�
�;�K&PR�8N8B�ϥ�aE�bъ �V\�� G��I�M����ŭo���1��6�{9\��9�$T�=o�$�'@6�
�E�+�C_��v��P@�Wδ��v���=m&�*��y����"C�Zk��+'�Nҏ�\b�X)���ǟ���Q#K��.V0gz�
���ȃ#f���n.P���S���V �=�;��3����h%��D��bq�Y��f����7��G2�����i�����I�Qsܝ��Ce"�>��h����_��tz�55F�y0~�t/5�dQL�f���\%�::c?	��G�F�������5�e~��l{�i]k�R�D�[�����8,h7�tҦ���d���n�}g�����?ў�oҰVc�T��pj������(��,
���5���,��y�� u��������/'k}�&fJ>��rŧk?�$*f�O�8���l*.V�-�"���x&!lSi���}5y��k��2�:��\�wT�3t� �_�ki3߁vè�x�Ŭu�W�������Z�r�C�nԯEt6��t�y��f?�d�Y���' ����Uow[E�dI����j��B9@`��
�-0TJ��8�8�f�p�<;;�S@2|��T������9Ro�T �_�@��C^�����H�H��k��xy���r��}K@$ә�k3�=?�|�@8�0��Z�f��cTFW�9��-/�k�A�}�x�i%��`š\(�(6��|�G̺�Wxy$��y�Z��Q򀰻I�t�K�Zۻql��:�7�M/�{en'jY����",[�,-=�׮	|	d@�LV#��z�!g��1p�ʽ�J/��NȦtP�C�Ki��6��!7�ĜE�Ϝ򞹢3���1,cXlxVHYEB    fa00    1880�
d�"�}�*>3�Ĵ"�g,�f.&'Y �P͆�`�ZC��.���tC���#�L�hUU�'Pn�À�/����C���,�t6��]/����v��lW�/���+�	�x�R���ɤ��]�q�S�\�4�>�	�^���yĦe��4kP6Y���gv:���9���w�֡onR�@����|����;.A�c�z��I�gr�e��$�C}'��`8�v�7[L�w�^��9��]:mD���H- !�J��9���7��S
�-�J6\ ���|��f�a崇k���]N��]l�b��_�m���3/n�:�YЕ�WF�xE��ދ�J)�N�
���eMc���_\5�\F
v��u�R����XhVfGQ=u8N|Q��٨�P
��(1w�f���fC�- X+#9$ʣ*����I-^q�d1b�	����e�`�1�B��獗ʴS���i��e��"�~�L�Ϭ�tz����N�)���*�.g:�mI��IW���^�I�9`���)s�(�-�q������ua߀�)�ߓ�L{���xZ>�i�a�Cbe�֋�/כ����z �\�v�K�!QC�nkT��v�o�z���e���i��v���KȎ�� �A`o�Ԅ����J>������Y��Nn_�6c�*�G�L���@f/�&Ԗ�ƳGQd2�3�{PM�8I�m{s/
/Q���{��HFr����-��RJ�{/��\aY���Mږ��f��烉�t��_�]Y-�\�p��S���"L�ՅB��=�	�e^����&�fn'�J���f�`��ley����>�)�����7��6*��v�b,�,Gd(J}�<B����	
Qb�Aٞ�{�����Q�\w�;�֋
���3���BCHC��N���3/p�~HB��o	&%�H��VQ"��aS��񯶤�o�^�\����c�t!&=m}H�����33��(���mV ���k��b��_L?�>��"��{�M!.�h-sd:����?B��h�ݽ#оj���5��2���4��E|�,��u������x!t��^����}cI����y����j>��jZ����*ݿ�7'N�џ�k�l��i�K�n�Nf�)�P���&����贔�b8��1Wfy���!��Yw�V�x�������Z*�e��J�yg�����R�d"G�Ѭ[�����^�E��FGt�a��oJB�ab���;����,��N�|�L۾K.���V+�n�)���F��xG��b� ϣ�ʁO�b,�8��O�1"�`�Pǉ��E-���|�[sS���'~�)�n,�&��&��f�T�j$ J��r���#En>��M�\t&� j������p�eLl�&�|;:8���z�GO�P�Z6N�@��,�r��*Hl�]�M�K� o
z[�{R�.�Gp�v���h�p��cJb�`,��|�@Q�P�	��[f}��]�>7��D�9�o=L+�h���W�<��������&����qBa͠U�q/���Y���:�^D�j�2��Sp�i�v�e�F�56\�h}o�"�zf�[p}2��w'_mKN�~�Y�tu��4V ��1���n!
;��(�y�W��;$�i�l.����y��X]�T��,��L�3��sa��J̹�8�lQ!E];��!Ӯk�*��� ]�	q��sh�`����ԻAnڎ��d���R��g�n�"
㓑i���k ��`I�n0�o�Gw]��%���Enc�����՛���E�yzi��#KKTc����qH�/4�����ږ+�6H�E�z�� i�,��Qd�0R����E�nr; m1�]���	�&`�U_��	��!���T�uA�S
LB<�/�O8�R0[�����K�iiI~)�1�0$�[E�z<=��ƌ��jA��v��&��D��am�~�T7��/:aML���cs���cU6��v�k�
s���Q,���<J>يq��{#{��r�ǅ[�|ꡏ)��S����M�=�g��z����G�m�^�{�~��:���7Ae��}�n{U�7:�����d�5"�{�0f�3�n�lP�KчH���W�i�p��!q��^�� M��ˋ�͸�މo[��l%u���V�q�G�A��*q����N�5��������>p�Z`>��`$-�0���}�Y�b�J����[�P�yfUxv8�?F/�������O��Q|�fX��b�s����������j���-	`�?�A7���f�����A�cP��!�:K*����  ǅ*g0��)�mI�	D��嫍&��o��<�3y.j�IT�3F˨��8Y�M�]u0��5-�����+D�e�!��RXw4�'�k�*�K-5�˯C�)�zd�g�����c�0{��^����N�OR	�0�oH\)�\<��%2����#D1}vy`C�G=�0A����Ն����J��yИA���g[0��σ˓���j�md^�d}K蟕�*�܊=�q�,�n8�;��mĄv��4�A��9���Ĺ����>�>�����	yՉ�2�
��4eT[�~r|"r	b�q�M��]��r���˴I6k��{y��Ep�c��<�ruh���҈�J/%V�ޤ}I�z���U/��yɜcoe	aEi���0�V����N+i�A�~%$��)�����a��&��D:m��hVx���a"� 
���H�G9�2��Rr�ikӮU����G���˺t�׳Q�{t5��v/�8�O���S��30K=վl�W�<�䝩.��G�յ柔��^)����#�S�[����S��M��ZVKZ��_�V(����J� �qOB�p_�;Eм����@G�{5l��5K��-2<��m�/p�Kط��
}AK� Ն ���x>�k[n�=��N��.���.���h$ǯ�t9J���Ex�rrwi�mxQ`��K��ݝm�0��L$B�Y��#p��M�xz��Y!
��� [>ӳ#G�a�"������i+��S/�l'�f�Ex�踯��-�%s]N���j���E�L��<UX"�M�8h�R��՟�&J���43�6JOn���l1����J_�_���c���1/6�Y,�*�q��ўB4�%��~�m����[ő~��Mwu-�ur�U�g������h�ͧ�:��|�%␉�o8�6Xר�3X��D��r|IW�5���R��s�a���M;��L\" Je���YH�(rG��'�	�N@[kVm��`X9%��-?[�YUF�5>j�1��<l�Y�]xNX�l��zP'�d\ػ\X%���ڿ�9��6�,�W� ���XnT<F��g6C�yF�[��b��:�C�l�$yS #��Cp\U�@��K�=U1�`w�Z�W�y�##b��ܪ�4R'Ʀ#��_��5���R/������d�_�E=�b����uu����nƕr����4��AE�?�_cT�ڽ\a�ij���A�^�%�U�V�"p7�8�
(�>��?��+���A<�q��Qdd�k����jU�B.Z_}���O�?Udps���]�>�˫.��I4 Q݅V�?O�� �ꈃ'���B��B�0q\�*��e�4�٣�'9p��;v�����C���g�4n���G���fDct|a�95�KBCn.Ѵ7NI�;���B1-�4�,��Y;#���ܘ��2B�ܼC)"�#�^e4Ʒ�ដ������=y�U�dܣ6$d!�ly;qa����%�-���[��R޲�)W�#�P��e��I����&�s��O��Vw,�������N��:M{���<$Dt�)�xdP��Q�����gVm�qmc�6AߪhB~����b/�ূ�k���27	!�����'�L�1wfsX�"쇶���㲈%폝���[�0�����<�����W��� hd|?ڰ=�!�抱y��R�P��S�`*� ��3HW�^�%�"�<̮�4��h6B���v3�['�S���.���C����K�4XX��G�x(=�M�>ʞ/y�����4'}; ��!R�F��U������yM&r^�nV6���E�$"% er3�+h��0�m+���Tz��0�Q{h3v��5�]��̀��{�@�f~���q��[��/���[e��ک��;�=B5GG�b{�6uz���q�`͍�����-�4 {lY m�MѴ��~+|�
����{��qз�4$Zy#ld��+�Ciи���}�nx&=]���'8���I帖�
T�W����m����9���wr�,�8��/�R¯Nn%G��\�ry_�]����x$O��>�*e*T}"�a�QL��	���+�M@𣫺���{t �������M:�\v&XR���:����#�[&hi��e��{�>�#�ce?Uw6%���*0��/C�v�1�^|-����E�VN�|�`+�k�MN%��yTat6J���kH_�J����"�Gd�~��)b	��Mk�]ӷ��(�eȠ'���k��IP�S���Cg�N>�k�A%'#MH����7D\Rs��u�����"&J�5��>6��H�P�	hm�0��3��2�- ���[�u�,���Or-4���y6H٪�R�Ǽ3���)YR����3tY��Xh.X���{!7�l���Y�Dx)
g��k��G�,~�'���c� Y��Ι'��F"z��Y�Q�CKm��I#2B�bh�����p����'?�K%���
r׵�ֹךh�x���An"�iPN)���Q*Y�
����BƩ�9~yK��O��-d�.��r�L���/̡:FF��*	��8��#��'�(rrv/|,ݳ�:��a�3X/���ձq��fA1��\J�	 ��g�v����"�j�~>� ����96���D��y�,A��٩{$vNX5h�o�7�x�M!���:�rV,�zɈW3�!�d��U��"��WBd��%�?i�PH*�	�j鲁����}W���q� V)m�o=�r�E��Y�
����� yB��:#0{�ڏ�k	�q�]��#W\*9�U���4�)s׉�O|Č`��]��lN�6�̌\ܸ\�b�[��1�[Ek�F��{`�������D�����XkLm=�Ul�]ۉ������8g����]t�J�J;{���A�`�!�sN�X�>��!��i��I���`���)��jS��}��O��� 8��iH�f߉L�Z�XxMy�4��	�PN��u�����ߩ�r��N9X�eN��x��m��3i4)��6�\h���!�������Z�N2�g�jx�� ���%s�����r�s������Ǽ��$�F��O_e�����#��x�G�m/���Ɓ�8_QedE��Z�P�O��]4���~v��x��&$�֍��~܆�G���پ*��N:��[T����*��;�
����_$Sm��b�e�s��͖`�vאaVO��"fZ��W8�����S��aV�5CU���*4�u�%��k�'�Dū3�K-��x�#"Sw�3���q�+D>�MZX�(�d]n�/�m�,}�+3��`Y�T�S�YNTm/�d������x'�x��U��"Ȯe�N����/�����?0M)f�=^f���`��Tc��M/Q�˿z%�7^���@�k�`�P��ͥ��Yzݶ�e��Pɒ�أ(�g���iiR�H,R�G����}KҘ��[6k��.6 <�����PPi��ud2�L.w�YM�^I/��&���z��گ�ܓ���Pt����\<��Ζj67�pb�i(�O=&�u�dJ>
��9I'`8{śM#�QƉ�^y��h�m�!*���m$_e0`Y5�]�K|/~�	���92I��}��J�ȥYp:��ۭ���ԯ�A�Ӭd\�ڷ$�D?3��^���q��?Y�>���������рW.u��M�Mvw���וb�ʄx^��4�%Q���a�σ��dlr]��k�N+��j6Q�s�Qʿ:T^Çe�`d��_�`�EN�?�H对��l�}��@�8�Ȼ�������S��řu� ���?- {��28<��*��$H�#VXx^F�=��i
��ӂ4�!���3���aEO&��iK'�2N��3��6+XlxVHYEB    fa00    1910�����$�s�8��Z�S�4u�$2���A��8D��e>>��ZdRD=����:�f�
�ܴW�Nޑ�f�l�j����7,�7?1�-�{�)QΕI��i�_s����#
8Z�LJ?�3T�DbT����C	 �c*3��ae�N��*X� ���g���������l,)��a.�_����Z���P`,��&�hY{�RdRt<�,��?��[b9����:%�=�������7�������>�*��;�5.ik��nQ��<S�lB@�aj	yP���Iu�\��ʥ�E�R��a´`s���������~���dpe)�
��

��Z�
<o�ѓ0GV��ۯWR�L4.Yo=�����E�C8m�)-�qь7��0�}`01���O՞�WE������Po�Կ��9:��72�Be�˳ǰ�8蔲��JB�� )l
��)�L�"R����c�ZJv7�8#�=^�«�uQ���9	��V��g��i��`P�hXV�BeS�b$~�q����9��w� -����k������9��h����s����E=�oU�/-:e�EDNx3���U�����GP��� ��Bн/'f.��	�!����B��t��d���C�&��p�D��́��~���T���+�]O�W�i��)KRSP�V�U���zP�СMNu,����(d���:#T�2�ۘ�%&���J%=3�a;��9D29Q ��p�J[Ak�Ff#�|"�aн>[G0��S�R�[:8���w¼[='�#���E�Պ!���_v�g��t���g+ ���fn�����0pY���?s�����d'�!d"�{��D���4�i���c�+d�	{�"*�����7��o.�Ĝ�o&��CNm��Um�D����~�I,�}�?� *(��5���!>K�?�O ���y��͵o`��Ԟ�i5+,H[�(f%.Qj�,��9�R���;3o7�<��?�%�'1��젚C���\9��E��e{���Y�1���������<֡���M���<�}�L"(�Rn�-��M�CAG�t���vb�T����b&�/��U[RS������ܳ	;��c��X�*o��d;�����~y�;��E%���_b���h_H�W��=��>��H�(���<���+ �!{��Hb<������+�*"l~v��(�F����F齃+�&phNͱ�E�]K��������_������tw�4bz���y����^6�	0�
jLʐ�����!g��u@_]��##41_�},0uU8Vۍ�5�Ҋ�g|���i(L�����1����ɜ`��O}qW �NW"kX�x�hAT���[b��J*���������1�]��.}a[�x 찷11�P��\,7�����P,������RIuC�U;�s��ؿm�`�0G�-TnK���M�;�ta�� �<��v���<Z�lpnQ��y�Ʌ�BF��RjpK���C�,���E�܍��Q���m�,)ט��f�-X��.��;����{�bt����B����!���d&������j��=�X��\lB7h$It����f�j�"9-9��&�ꇹH��c�]�lWd�^@n)j���tc��!2^%�&�6}8A�<Џ0a�5��+	~�W�&э�7%ҟk��,�n<"�12"1�!�����J�4�ĮM���Oj+N}��ɪ��8I�v�s�B�E1���:u���۳�Fې���=8+5-�5�K*E�xRPj��~L8��5���盇�Ϊ�(iwL�K/3��^�>:�5A-X�iF�+f��HD$
��>N���y�j����?i��:-x+�M�\Q#S.��`��E����b+��6�:�H��źAI|���B��e���W�f��HH��R�IB�?��܉�/?
e���C �;؊ש���F��7�cW0Gt�x�"�����R^"��G���Aʐ��WE�V;�쎺��S�O�U�A��0>܉,g(�[`��-僕�����-u�̍$��� ��0��>�3iI)?@���`sѥg�R�M��+�=����7�0��u��|��jʲ��Sa�g_��\_���9 if(�ªq
��x��U��oy?; �L��-A��*��mn*�X�d��r��T��H�'s�dG�z[v2���t�7�j������-��]�F36Ie�
� �Dj0?e�d��x�ͳ�^G0B5��T��f��'��|�QɄ4P�g	�π��ӌ�s���՝4����^�:���\2��%X��Ƃ��Qj
G��]�̒v��I�P,��!h�7�A����� �s�p�^J��wY垅��y��5�:Ne7��	�s�nz��/}�ە,EG�����M��5��D�	��(��XK\/�z�,�Tk����A�߃\:�q�q��B�����Kv��`�Q�1\'!�}�c���}
����'�Ң��L9�MbR_a��-4!���r�Z���vQꨠ�2��Z �c4�*�<xf�������aŕ.�F��
�7%[yh��oiI�!�-�t��כ�9�Pn����!��s)�%�)Ƨ�׍��tg�Tmߡ��	&^骝��h]�i&1�FT�uK6��������9�����9��%�~R!qѕ�����g@�b�tC����ƒ&�;@��iC������nH^�q&y�N�CmgZ����@�G*
�E��ὓ�َP8DoVR��>H*��a=3F{u;��@��u�؊�+Wy&;�79��^��E�30<(���2��Q����h��h��As�K�G�T�����(��ߨ�q�NH����f�q5�q�KF�����;�PY�~F?s�{
ϯ@֏x�z��>��%5_Ob�3�7nY:XV������w? �0e���+��w�~F���� 
Wv�.��$��04n�������-霸�]і*�����,�;�#���*l�9�m���j]D�P>�"���D~v��͵XǕ�^�de|A��^�\��Cz��P�T&1�Mx���3�o�^����)�h�4�5�]w��îѕ�P$�yA�I�~�=C\MAN��亚��AX���
�B�q�!Y��2�����z�O�d� mL�Ԣ@ �SaB�2(!$��!�yX��JJ�xU����&�^ˣe۷�y���=��[C�j�3�u���</�h03ZJ�W��XS	�m��t�\���L��s�Q`(z����f>(�Cw2�w���>ZS8F��"z���3~��m�V��GW�%i��b
V&�_��\��G1��zv)@jr��F�K�����V0-��Fb ��QN[�e�`9&��e��p��X�g��H����$Er� d+3-�AfY��w��k��>�~m�=�cw��Vu���w�z|�O
C�?�t��)�`J�^��͈�Ѓ�Bk�B1����}M��� ���`��F�z`aҤ��Oҗ�z�=�[�2�B}��5���bOS��Y2�H/>���}X ����GͮQe� I�Z�=���1�P�E� s��Чɖ��rt�eT��p�|�,7p�a�1Fa�i�2@.DH�D�1�'�Z��c6�W�A�~n)Q�8�כ�g't�y8��7>���[���Ĕ0g � ����Z�;\?\!�؍�Q�Iq�ݽV�^��_�X�s���yr!�#<�&��V����Lc 3F�[��� 6��s�ڵ r[���(��:�n �Ū��j
}5Ŏ���J]���LM�Z�c����IY�X�g,c�a9 s\%��ğ�����4%�V��\j�?���v��;Q�}%(�8q�_�ᭆ��©�h4(�x(���Y��X��	�/w�Z��=����d�=1�l������!��=���7(y�l�X�52�R���lU�g�TЙ^�w+(�*��d������qZ�J��m��wqR��JT��/-�����T��gI(E0���)�+7HFh�g:t�����s��䖫��J�u �ǃ��EO���A^����|&��=���E����H�t�����M�@��|�ٿ�!�O��8�Z��T�ד|�o5��v�<�_������Y�,�<�bzi�n�I�H!<Y�k3�n=��u����WOy�z<�'�H p�]2H�3k��_|	��w
썩�������tKvP��"���HSGJO )A��/��,��� ��J�^�����<P��𷟗4�/̳�1l�z�S�ɯ('n��H�Mn��l!��W�eN��B�أ�q�gY���.<#!��1�dm!?�A~�δIb,�g;���5x�f�p+c%*��
����8>�D��>�7w�f{�쿹�:���&�I[A:� 3H]��b|�w����
�*P�+��A��O^�m��K'�wj S7 =D��m�[V�����!�bX� %��Y�����J���B�6���Y�,n�:HL	u4�vaU�<���A0���D�?�����VB��(�ׇ[�^1�D^�۽�u��S�
��s�-X���|ݽ��+\2�Zr�w^��j�z������h>C�J�ޢ1�9Z9���u �*��yP�,�!���"��˅�:[3�"5��7����]H��U�i�oj��#��7R�1tCA��?VDie��TW�'�ݬ�<8Ⰷ���9��h/?u�����'+��7���.�M�N��_���/κ�S�J���:5i�%���4��W��b�N?����&1�\,W9�	=�D螚����D���
����8� ����J�S��!"밁]eo1~�1�}v�~�m�Q0����CF�:�@ᤱ3�"�/�%�ĉ%РH` ���)J�]�&�c��9�����_Q��ސ����elaUw�.6��7��W-�ck�S��X0��>p�i���8�;�) M���DR�f-��0d��u���(>R�^P�o|�u�L���Ώ�춰D�Bي/<�ߊ��G嘫gjK <����"H`"+�׷;��K��� mU��������.iN�����1���o���xO_�F��zy�;���M��GSDe���5��G�5si���!8�3���|�U~4"u�s������iݿ�&�q�-S��F��t�XOj�6�+`!8���_�x��Ҳꓟ�(G�y�VcP}�>�
��.�,g�x�y%�nR���8T𢅆�%�؄��	�0�a���z����N
�
��r5�ЇH����k��y�(#9��cMq��.�i��F��`a$oA����~Ÿ|��e��:#�ˤ�TC��&��k��)�e��·њb�G�x�*�iTlcQ~��*���HЬ%��g�o�aغ�C�@[;��B3�&Y�� ���]J<Ȫֹ�2���8	rx�9D�;扝�X'��ʽY��^q��ݝr��b��SϜĄ�Z+Q�d;>�6&D���#�v��prA����=�4�#F�.MC"��=�5rcx�|�m1�ߐ�"Fc7j�RQDZP-J)�c�~v7p��O�v�J�qi��(�l��dY�I	P�s�ʀ�o$������04�_Q��Vf�+}���R(��4����8'��M��FDk �=�ڃnf��7�߾�s	|��D�] ^���;Z��}t�TO�����1�^F�����LJt���v93f��s�)��a��/+I*���sR�;�
�89睅�u�G�~Z�_��;җ���Kы��bQ��$���z��בa'���#��<�`V7�ˇMM��?��LzB��ܒ�-;�7fK�a�)!E/��-C��@���^d����@����,����P)7�չLQ���'93��c���)Q��Z��򟶦��܅x^M��4hb֯P
 	׾P>ַ��Ĺ<k�j5v�CGޒ��:ڮ�ٌ��G}�"ʾ��(�6Q�����_�9�/+�Ġ2�U$��&��˼�f_l�D��F���=��@���B)`���BU0����NN�Z����c�\}�_r�?�=�36$T�E�1�Ki����@� �]o�6��<궴���\B�YϚ�@&U&`Rr��˴�5��~M��$�m=�`&��c{��	1c}�� t���X�D��l��T�֥��5�a��#�y�V`�u@������YlE�2޳��i)\ԖA��[�9�l�?�c������7C� �����G6�5IB���!��"��qx��SE̵�5��5!��9�gߊ	�꺓m����b�~�D��;�>XQ�	:��>�#W �g��WaH-�]�@�P.F�"D3�e�
��'��;�o���BGl����0wEƒ+P�S�8�- W��eT�^�XlxVHYEB    fa00    10e0�1��|�����̙�;�F�ܵ���������ݹ'�$�b��2����/B�4�/^-3��h��:����(!�a-�8ng>�"���Q#�^���!�8���M+�$`�և��d�}�=ʂp�K��Jt�q� �B#D��1�)	����ԕ��ᕯ��L���oT�g��iQ�������3G��d4"ǰM�S@E��~'���Y��)J��ā�.l�����G�\�����	�R��&ɇ-U�F�}.����H]�d]j��?�G(��ek+�+tm%����1w�6!'�l}�D�y�[�O+�;���ʣC'�;%��/oY#��v��Q�I%�Ml��+�YMM롚x%��eS׾k�T�;x3�}2�6%<W��
0I����}戯G�=�Cޟw����3�*q S��Q�����Cp�P4-�)�����H�|J1ܣ�ߛ�~������q}31n��F���,��U96�Ɨ�bI����Z|��+�J�G�r�ͤ8ߏ�s�6�qH_�
�5E�.�АnC�)�����l�T|Z��E�����?�����yJ>y��p
���L8�qf�PЕ��;D��@�]n3��&��=�Y����6�փ�}?OU�����A~X���S
n�x3�F����ݨ{3�_lॼ�	Y�uwn�.�߹e6�j압fD�=޷[��ފ��^<-qxE)�����F��Ĝo�q��̴FJ$-rc�17���.�l~Uj~���I�y��x��0,>���TK��srqm�2Ѐ���n���p�z����Z!��[3�K��چ*���Pr�
H-r<)V dw���ҝ�q��v���VGzE�����
��|�	�k;��E��W���
eѸx�7$u�O ������Qh�Y&���lSw}|��	�j��[��;O�x�i4�S�����$�3����:�����Q"���	�E��Ec+@@">�d&��$�ۛ����)�F%����/�gq�H��ͽ:0�N�SZ��ߚ$�*=����5�Y�0@͉��K�B\�uX{�(��g"Q��]������,k+�)s_:-�o�~���$"3�oJ~D��!�oM� Z�5������P��|����"b�"�8c���&��8�5�"��������[�V���"�]P���yMpq3���/�����үc�.��?E]Q��ۣ�z���`�ā$�(`'�Ã	.�#��9���C�N<��Y�Y�
��lcT4B�`�-9f���Ǎ9�Dm��<F��l?�֎��i�Tx\����7l��f������$I>{D�r���pm�R�;`�����1��;a�z�N�@�	�F�n���e�>^\�`�8��S!Ы��h�|�_2��D��B����$���!���V߸�W�Pab�� ~�5������:Me��y���3�ٴ7�2Da��؇�a/��
�G�$8��?�/��ޑ�8!��f���?�ؖQs���l|!
�7�hǬ��������hq�Õ`t�S�;Sٗ�B�"����v�fyĵC�p�?�|�6A!��G�k��Q�Qg ���W� ���T(Nu�o��;�NsHT �w����.���a�򆀝���b����+p�<��Ҭ�zY�+�L^�J/.(Et�JDI�UA�"�
�sє!��^ьW3�l����)�#Pnd��KzIR��,��,� ����4LG$���Ӥ����(������q:*��o���j�q)���%7m��ۦ-)w�)9l��ʸ��C�D����cU`�P����i�H& ]h��r��+�܉��Pk���I=��*���+����T㢫���7�x% �{a����ZdL���Q��o�8:���H�<xBV5�[�m���X>�Wet\T��}~���sjV(~B7���W#����O�(��qꜤv=
�mD�MhO��2t�s4=ƳL'�� 4FB�pM?V�5n�0�2��԰q�|��:>�R��\�M����3��F�
��__�>�b�o�כ����H%��pS���Ԧ� ����̓`�[jT]�>����0���!jc�6D��3<�~��͔�+�%��}�F��(��E���|�V������!�чRQhs��\�TLȰ�)b7`�_�@ΜU��/�<	����ϲeESM�x�����'�lN9n�v��O�eH�8!g���mm���Ꭲ����Cp2����d�C??�Sӆ�Y��A��C�H{pΤ���b�4U&�ůd����j��Ï�A���\��>�ǔZ4�6�G�Z��#���
���y�Ѕ���l�S�d�vJ���$C:�
V���N�c	�O��K�y�p(��o�~�NX�I?��
֕��Yeg6��F�c,�,rN(�0�����pdX��DK��$i	�t�>9��To{(�z�:7d���,/,�$�!?t�&(	�v�]���`�����)��H^�͟�s�����۸��4R�)-��Gb�̵ʵ1��{[�cx���i��G����U�;�/56�=G`��H>����cA�2��J��X�B�B��=��D�N�)鮛��'Ӱ�W�7�VF�XV^Δ�+��t�b���~�wv���,�G�4{�b͌@�L����l��c���	y� ��N;��A�,�yd�V`�x��X#Sb.��g�b�{Rm��'����@?<C69�p� �A��M�# �Y#!��+�wF��X'�:$��|�R(�+�1�?�����Qsl�+Ic��̭&j�3�P�|y�F��	IhL-����e9�ȥ�^�d�4R�D�)p̀�S�A7�v��i,�/�áLi�uz��n>�Ţe��3����ױll�a��a�s2�!i�.6? �Q-��jW�1���[%�"�*���D:�膮ˇ�GgՖ�^���Re��g k^9*K��|l��3m�7
�j�C��`�"�ԟ�7�E�q��w�n��YO��8UY�`#�6��9��嵝���݆$tݸ�@�ӫ��<�!�*�J\S�p�ir��T�@����Z��P���	Lbv!�a��h��G��<�&9�ܖo\?#��D�D;�Z>{��� 4.N����
��%�t�#��ڜ���H=p���{��pE��Y#O�&y]~��]��2���&�h��H��=Z�",[��2�%T���↳���cPZZ�i�I�d"����sw�vOB�&�f�lq�9g}�A�z1���������JQ����Q��M��A��8Ӭ�Ɓ�"��V���ȃ�&%&���;�"�5|��d<m|����5f�'^�1��&')��.@�Y)�Bp�A�"{k�/�qѦ¿Ѱ�Ӱ�$�T��ҭ�S{�sS�u�L�H?V}�t	��X"�/�[�ȾꨂÍ)��=O�2�[ߕ�C�VW����=`�y�6'��gDx<���m毬9ә��Hߍ�D�30�l������E_�gFr2\��i�O�;w�C����yqmu
i��UIN�7�Mz�{$�o��s��M��gbQē���q��w�<$nK�a1�}P ��gG�]�Yss^װ���9�i���t�����f6��'r���w�I���!�e�_���8r�Չ��b*	�$��X%��)����Q����0�!�'�n[����@��@O�o��h���E:�`��R4T����{&4"2�+Y$��Y9�RP)�CJQ��C?h_U�%Nkj��
^�ݴ󆃻�C����X�d���J`�p%�X�DT�َ"w�+�V-2��b�6���߸`�Z��m8�5��|�4��аa-9DE�2A���݃�y���"�^^lKbo'�X���U�A9Ԓ	��ى���"��1ۗ�c1��7�����ms�6:�T���5en�'U0�j���g��|�^FԳC��G�Cq��d�;M\��,���ᗀ�>�G�=��I��KפE�~�7�#rn���#�Nq����&J�B����Lb��=yp\��T�5�����kd�7��
/��X��<����>n����N��(�HΣX�"I�0J Ë������8Nc�yj�,�0�f��5�ޠ�p4xe���bf4!�G�a�p����$�@�k5�<��v��Q��k��@+vz�N�^:E��垀�O�48��?� x�q�s[`��e��B�@ԇ��>7m�O��<ڙ��$=̉��<B�z�p����q5�3S�j��7>�L�&=�'k�r�gE�!.�Ro���_XlxVHYEB    fa00    1860� �t�kO�T�,Bؕ�O�P_��9��O���m^�R"Ҙ,X�*�R=�1�*w�9�	��O?�	Jm��|����z\[-JzO�)��e��f�7N	E�_LȲE��5P*�]CL��f%�;?|<�=<T&��呦'ӱ)t3"���zG�,#��!+�a���y�j(f��sĉB�*�'dLT�C�C�T� ���8�M�l�&���i�IVѨLF�s?2%,�p]/�LF\��!r|� ��2��.�����yj�MyV�Pqn<�f���©'V9�$�f3on�8�Bj_�%?��4�iH�8W���E��L����f2�U���eb� "���v��l�gT�����ޔ3D-�J+K�����qh�|`o�v �+Yg�GGb�A�󆉬	��Ǘ�:��_+�6����X_J<��5,M��>f�<@��e+�� ��I�D�d�M4)��e���Eq���E�co	���ʷ���SǐJ��}`mn��Wr=��x@��^��1Tu�zWQ)K���!o��*�X��n撞�� |����
(�b��v�����J_1Q��>7+P���KPh��LAE���X[�׺�.�)W�5���MkV��k{�Az�����n�*�����#�c'棙m�gy�V3ͼ���k�d��e��L��LYg�����?�D��`��m���xB9[ ��NQ>�`���R�|t���Ю�/_вؔ�oi؟����T��|�?�\��]1+�We-h��dq�-ѩ����i��ԋ�}g)>#�'w6�������N��+8�Iق#��O����\�$q/_�]ll#����.�B�H�*��H�%���h>������輚��V�}�����PZ���I�a�?Y�q�Nq^��f���+��,�`3���Ա�F*���z$��[Gi��	%3��=AGE)�~!Y��\I�k8��*�^�|�o~�nr���):3B���˲��4� �/�$���`��!��ݍn�П/����2g�`�8;//(6�<�8�)��V�9LvC]��Յ.'�|������M)�����mGP��d4��:�v9_�y�
���K�a������!֋Mb�#�	3��7��suW��p�E�L�tc��N�|�(r��t^�Ƽ�sQ�*�K��K���hlMz�nu�Alw�a��u�n�M��9°�n�zD2� �0ADRn����q����+�i)�����i�_�`�z	T���žQt�K�6R/d������;	6�)@ߜY(��0���6��W��r�7	������\�2Y>���,������3y��T��u��U4��o�u_E[�=�z�rf�pct���Q=�I�I��7[�d�˦�HNӐ>�b��xy�=��[Q�3*�A�+�N�Y��;�U����ͫ ���(�D�������"�߿hM	?�֝<�ÅU��ޔ�%֕�*���Ԓp�L���Lhp�/5���L=�Ƭ�4�zR���Y?_+��@���H�Ϟ ϟ��fN�F��;;%�naA<�:ќkS-:��g����M��]]�|L�v~��늮uL�$�[m�G��r��&��h��
&�-��Ɯ(�~����y�Q�P,O�e/��V�<"����=xj�A~p[x�3� �����v�`�u<al,ʹ�ʩ�W�Q<=^���� 5��ƹF�?�ˢ��N}��9�<���'"��z����;�<oO�<�,͋�
S^�M�jD�p�A����1�>r^�$U�l<�k�0��j�&<�����J��Սu�*����ϯ�cndr}m(&�Ō�0�����*G��ʔ��a���b=���*~�\�h���6Q���?NI�GEU�O�f�A*N�G�%2��"����&pTvI�"�f��Gˈ�U���BT�ޟ���hC��l� ��ZV��*�4�l�l n�q*-K��:9���훚6��`�YпzC\��o|"��K�ñ*�=����s7�O/��R,2����m	��,[�Eݣ��^�х�d(�f����5�H����N	B��,P����p,���9�9 ��vG:D��]n�d�J
}�������q#�g�/  ٝ]�u��khx�՟Z"�<~�:�\�4X؈�/vX�y`v�6\4�Q�� ������:�����g0m�>!��e�Д̊z��N�d�J�0ޢ�����6U�6hh�#qx�7���8g����Ƨ�1/h#�3�.	��p�A���Jy]���J��/�J�α �J�"*EXsگ�/���W%�5�D)�>ɳ�G��N�A��C]�e��5��Q��F��|�M84��D��<�U��Ճ��]a%u�f�T�'�!��Y��������>!��?�n��~��0� �k�}��C�7�����>X�u�F����ZMX�d[��B2��y���7�����6 �tF	2<ۢ�V�%�DL=|?��-V�r3`!F��[��&��]�i�K�40�B�(�?��ֹ]��x��2߰�U�@m �T���u��$���`����# -�	��*�U�+!!��m��5�$�����Γ{��?� �3���z����)��3b��̦f�x)@�ƍ~��>k^ĪH�>NL-�m��z��2��v����iC�z��8�b1���b��oڠ=��v� ��_Vم��\�3�P�I�U��4��P1=��$�X��XYc[� �/���l��j<�?��x)����v�:^	�1Q���n�x����^j!�5�)����+2b��_҈2����s�ƿ�R��_��k,a���M��� ��o��[%���\��*�ڋ���_ꀍ��`�+zZL�	���7��G��Y�Z���g��qV>�YP��J����/�LbO\���!�(M��9�a]6�"+�&�ItRk�!�'+�ӌڢ%��|N��g���ѹKͷ�� ����\^��U�X���� �����w�J�I_F��� <1(^�� ������:����_��{�B��t���S'�@�����u��Q��w�b�M�o�� 3]S�Uq�g��W���������VL;&1/9p����j�R�NW6S���ōF>t�����ϣGʍ� +���!ߙĠn3�CϜ<�)%9:�TM$�;�L�X?�2�<P�~#M0�#��c
K�S���!⾉���a��So���83�7���a���S��s��s��#�OTa�x{���F�l�����U�m�*���!��"��`����A;O;Weui<��]7���R<6'2�R��5��K��iKo���� ���ɻ��ğ���>�f�=\���5G,���[,�.������˩��p[���{��q`�Uн�������fh3�}�c�^;�7��h+�V�� �3��RU�(��I�.@N�H c\S4#&9G��H�Ӭ�UߙoBJ+�z231tE��c&%�}���1�mnҼ3	��-������i��N]�Q�Pd;6�W��TAPc�lM���-�0I-���<;p�����{ׇ�˗�Ϫ$e&ʫN����R�*49�����o
E!�:Q-���V3�F ,�1�{��'eK/��_:qA�m���k�8L�޻��ʸHn3��H8�~�? �SU��o���~� �n^��;h]ޒ��}�g�Kï�Ё=Jn�V�h:��pf��e�[�%H×6�0:�������/%)󔻽88
0L��Ξ�V�D˾� K_��S(���)H�-���xk�B���h"�`�P�{�d���_�yS*�Bכt��/m՞y���$<4�e�/��j����R����N���m����V�^-�"����}�^� ��K
�V�L�C�9m\�o)A��-�S�?��(%~U�T>��9��*��˨M�H/��ǟ�P�������η������[��q��1?t�+� A��\�+���ƫMJ��J�g8�p�۩���x�I�BP�Cb((���'�2|�x`Sl��?�1� W?Co���{����+T���N��Y�aƲ��л��\"0g�nݭyj�D��qٗ�z-&wc&Ta{��O�K�H8�<Rf�S�3�힤7S�{���s��4��!64����3H�s�����M�2��80�NSU�N:����'8�@u��'�KG�8��C�WV5v���7�@��<��.���=h���#E��쓰g�Px�_��>4�o�i�4(��C�Đ�}LXJ�ڨ�!�_:M��N�>0K�
��h]��"Y q��:�ͻ�G�h�E:�J߫�G�[�9�E�q�������nj�~sשI��t�"�ߎ1��!��ިi��iÿd�>S�4]c?�w�D��mZ=����-k�;|\�O���(��w��nP���@j�y;�
r1Fe���C�Ɏ�?��9����U7O~����8������(3v��|С ���W�%�ۜ���Q�[�ug1/����K7׹Xٟ�ᆣ.����k������h�9�-���\eBMGbvG�3V��ͷM�"�mNj"ʳPŻ��������*��*7<��5=�����d�s��Dĭ�~*���>2�%Q�V
O�\K3)����h���Jtl7.?��t
�M@c�tJ���9�R�B)k��{�2�����uz\�HbB5�At1��bs����m2W� �p��M11��)"�J�=�e�3c��B�;͢.�F� TK�+\��ڼ���{e�v ��1z"�A+&�_���� KÜ}��c�������5>r��Bnu}C�Óy�FěU"|�D3�@]Cuq~���fg����-�8 i�.D�b��]A�`t��}��nS�:E��H��'�J�Ic�2Z�e���'8_ ����Z���G?x��^Nu���<v����h���ֻ
�_��7l�|�"p�R�* �1��p�7N�]���E�L�Gs��5+=�l{��,��Qm�-ۃ�h9�	������\ŵ~�=
))l���"�b�UM�73�Ͳ{>����7 ���o��+�݌V@���u�L�v�0d���U=��+���I�S6__p���'*c���E�6��u����0��ψ[6��[v��$�JJ�ƓD0uA�Uza}zxT�\� �cM���6��D�8�x�Bf���R"�xi�y�f�iZ�E�l�&W����XW��|X`Ra�;�!��d�MN��JMѽt�ӫ��#�4"��FF�E�E˶R�V��z�:$�v����g���(?�%ns��mU	r��J���kw�a@��pA�a�/G����v�dv�U'��r�D�ʣ�@�4�\fq@��e�b��k���'s@���V���FNy��|���6�c/BZ+'̭��A�p�����f�>B
E��1��T��Q�B�{uħ��,V��n����@|�Wr�iM���6 E����i8�/Ydm:ɂ���rv}� t��,cS#&6��]����<��@ǌ�l(#W�4(�6��ʊ#I���<|e����M���(�ٷm��n>�Ԓ:n����� �J�I��?�t�xy�mi"��ߪ��nP*�wYsYF�sXY��y�;.Ծ����-�c��ź����1�L�f���9���}�*�Tc�̴n� ��k�O5�"���CR;��l��|ȃ\�Gm����%����z]��Y4��� ��u��.�L|w�֞�F�D���X�pi�X��t`>N:��-S@~�c@�`s��i�˓� �W���p����"�)��:��A�sI=}��(y�z��L�{��Ӄy�:��s�p��@���a��Z�G^L�D��r����ĺ���Y��ڊ0I0�S�@<:TJJb\7�۴E�'�SD��{��R?���U�@�B�şpy�h�u�WB��X�-8G�����I�-D�����X8�X7��-�'���ʿ����u�d�IFҭ�A|c��}E��É���ϟ
_�9"�
���h�F��rl�D��p��D&���I�n���3� �! Ĝ��W�ͣ(��a!EM|^�.��.z:�,#��FU����#~߄?�-����a�I�1���Ѭ�s��붴���b����~��?K���Rz�j�u�ٳn^�Ӂ�P�	/��3W���XlxVHYEB    fa00    1720���p�Ʌ�b5<�<��12�m�#�!�~k��N� ����
�YQ�a��z�|�C+:�8��9��aV%��:nE���E_�Aq��+8����:�{G�E	�\���}{M5������ �v�[�>w�xW6�J����tԊl=���Ӏ�Ŀ[_����S&�$6�*��s[6�#�^\�{ )�}j����}ӯz��Z)JQop������_�v�F-gn'�W=���$���;Hl
���y��e(�d��E�oD��3�ޏ��6�B^E��/AOt��g�5�����%A50�����=��#�9��ٛ�ujTTԥ]�)ҫ'#w�-g�M��ϳ�;��v렆�ja�r &_dAbr�Y��_���lVyҚ��y�<$ɖ;�q5���ܳ��3iF#����M�O9OR4J�����՗�
���"Q0�*�˱ca��e}��Ӕ&g��D�d�d�#a�"�\$�����bH��it��>��G�I�ק{��ҁM��N������,@�ST���vf�y�%|�*<c`m+}�|�6���>�H{��*�_�\;�ڽI�#9��������eb}���@h �3`++Rh���έ6�3�^����;�-�_��.2�\4�:�q��l��pP[	 -p�HJ#��Ք�n�{Ug���66hʰ��D4�i=�?�TߥB=�tv��f��x#��!���?�׿�����KH�=����u\�.@�ῳ�dE�bE��ț���,_0��,9�'��/��W��&�T�@rA�4��f���ꃎ�d^�L0�� [�@�]k��R��|�q���s�����U�ሔ4��$l�����kL��U�g���Wq�����!z�ՁZBPR$pT?	_���|�҈oG��L]u�k�j��Z(�ߪ4� ����}��\.&�?���}�-&/��O�m�Q��ܐPP���M#q�	�M�]��W]D0�n?S��ꛋՄ�h��b�:���f 6���]�.M� Pȅm�
�<t|�H~�?^o��隑aU��S'�0(g�Ou���`-�fZr`%�np�+"a��x�G@�G������yp+|{�9"���>ޤ�J�\��F�BN@ٴpV�����Vr�L����cD�ޡ�:�FعL]֧�O-Q�*l��m��~�E\'� �s/����F9�aM�(��x|�RQ��8;��x��|el�A��͕mm�y�0?d@���eL9ۦ��,���3;�'|�@�-.1��ǒ���g�
�����W�U7����A!fr�kVjGr�%���.c���ƪ�,�XG�3��1�.(�f�K�g���Sh��D�	\�mmә�i�=�i?��d�蘒<]�o�fp���R1Fo#hmx��yr��kKl��������ڔ��79}�q&H|4ß���soM������_�������b�*#ZR%���� Í�	��0����t�6т��a��ԟ��#o˹�T2�[�K��V�_.�t۳�]�r�d�d��j�D|[���d#��8r��ђ�v������#����#�̂��DYܔvX�]|sq<�ڬi�Nm�����([�����U�ƞ!��.�fj�a;3S��ܼD�F��Ԩ���w�3���	���H��r�-A����n�o��%u�J�V��[�G�/����?\	�p��%�[�7)!�!$zp%���`#�4/���`����l�^��!��*�*�����uli7�d�+��O�
�K��s�<��0"i�YK0��ީ�f&��y����?P Mp�`�~HJ&��l�CmE�����򗐽3Mv�0����Stv�m\��M�'
�01霶�5��T�	r��A�ʂƚ!�]$��T֑�J���p���[&�\��[zKbr���/L�M|��;Ao�+f z�ޥ��\7�I��+��8��M[�^�ܱ�-�v6m��l~q-�����b��t�Y��]n"�v�y����xL�N5ڹ�����P＆�~�A҂��;FX��~g�Lo<u��EdUb��1&ػ�λ=zA�.���a��-u3�bq8�;���({HEM	��"2�u���������@�ƾz6-��MB�#���_��iF咜�҉@��d�ԗ	M�WfO�pr�dA]C�C��.�))��%�v�뗨4M%�e#S}��o&Y1����r�vI�LTw	x�F�S*4�oY��/`��=>#��q�[U��{��B�|�:�YV�h4<O�$t8Y��k:���
�#>hOT�������^X2�-��nqg��t(��gi?�h3�+j'�M��(�eh��SV�����nȈ��zu���+�bB�f;�j�bAR��ےݲ��/X��k�����;鯼O�~-�Xc��щ��g�]`��.b��x��7e�v�vD.�r'h����H7;�~/UN��3R�Q�^4�y�Ny~$�K�	�!xƮNB�%~!�۶�ic�m�fR{��ό�
����m=�6�T�M�I�®�s�`��+8�ս��X]yE�Y�D�@Ým0LvB�Z4�Ad���js>�Y���CW�4�j�S�AjEK^�!���|�5�4@Zm&P��Ib�W������]H=�����Xwl8]����ԧOT@G�Z#�٢e�E����#S��N�r�a8Ia����r>�娛O1ܓ�"����El`�'9�ߘ���p�z�U5B�=�o�ޅ"�! �j�l����L��H��(��T��H�|$��P�O��	Lp�s�,��lg�RS�<g�R"��}�ձ��qd��x���	�����+m_q�ǹl +�sv���'EIG/
=o�xq���Ɏ�_�S� ���范��s��d��x&p��%�u��h�������a�ŝ`߿�[L�|��.�m��`��'�f��^S<t>�xq�;	Ax8��Ғ�#��i�iu���Ι�?n*<A�{3����+;�S�3,�����͑R��pV�=���ԠZq����{ۉ{<�'�K�"�B����{`Z�pf~�t��rJ}�TY�s�Y�7�C#���6�"��F�F���U�R�C?zu0:k���cH���H�ƃ$ f,�����D�E�^���|�:�xx�$��>E��9�֭� ����HK	S�҈��{G� ��HO~6~��DP���N�1t�2�"o��=f������%˧�HG����`�7�V��7�wJy)��P*R�::Ў��&R#4T�5���̒C�ݱFc4��>y�G�ë���jF��9Pm:����u�g!�8iǙ�nx�x�T�VM��E}3���n8�o+Q�9��\=MX�Lɠ�&�m�͹'�\�s;Wf�p��k�
�8��`Ό4����X3 ��aX�P^)��j�-����b����m�vђ z���޶�������<�}ߖM"<Qmھr��/?�;�}qw8������"���^1�j`���������G	�F��s�Ќ��<�+�]��"t̻�[���Lp7� �]���3��V�������mi�CIGHiWuWE��w�ñ��9��x^�.��j�f�C�*���l[�&�-�_�a�9#���x���H��h2�v2�I�Oc�h��5(��!��8}��B���ݥP�Uq��Xdt-���)6p��`z�| /���X㜘{��S�Â�s�x�l�.2�֬� �+ra��Md��m���V.�XQ&{P�z��%?a��U.��s��~䴠�.�祍�{A��d# ��{5�  ��bC7"r�f��,r���
�%���8���n �Lr5�5���72�0�����Vw�~����0�^��2A��+䮎y�����\����&&lOA�iW`�րw_z������`x�L�%������cRI�����8�k8� |t���ż�u�\�~5��K��Ո�}�ui�z\�X*�iTe��LE_˷FsL��#��������ܓ���TB����^^��N�-xj�]r�~
u�ɿC�v��o ��������T�,�U�vz����e�̪�K�4=�[e\�Z#@D��wTFb��6�w�rw��ԛo���M� ���N0���*�MF�k��NM���Ƃ'��-,���##b�1C���9c�
�~�I�Nq�fqA�Ԣ�:�wp�I��nb��Nh���A�<��p���Wy���k�%A�m[xC�L6���G�"���r���@�Q@O�nȟܖn�v4�����U	g(��'����;�l#Q�{햷��Mc,e��t$��Q�'��ޙ~"����@M��"��(��ٗ��x�+�}{����@�;�Jƚ�J!�MO���>d>q���&@���@� Q�]몾�_�c]��`�fm/u �O�:�K�['�K�=Qu�&n)f:���|�}<}{����^ƃg][��y
�Ŀ��$t���?FI�o�-��A�Ѣ}\�¹�&]��@'Sf�oC�W��\0�#E���!_�ݻ�2DU�z���@Y0�����2bEBK� ���/רN7��l
��2�-�	m����
��m�ᾶ��m,�)kIQ��8d@'	���TcM���N�o�Ԅ�q����ǹ_2N)����V�W��ƴ��
�SUDjS�B�`��9�H��c����GL��(6� P�#~3�D>�3=�˔JIF�uC�Ȣ��u����g�N\�!�IU(o�ۅ��J\�����a$��Xܬ}�";�pX
�j��gt����f����a%D�o��X%/�'�����Y;��>5��#��*�b������G��v�K���Fd����)��P������������hWf��ƹ�x_�'=Uҏ}�U�����w���b�Ox�,y��~Qf�L1��D$C[�:e8.���TW~A��o�p�Š��]\-I~�t�ȝ����p�������*�����`�.0d��
�.��T����Im�ܶG,������k0��}�	�;[��w�EFӝ�G�zĸ7�y�����5:�C�=*�V�+�f�%b��V���]��bk�U�_��64��3ʯp�i$ߎ��1H�}��?CL����ʵݩ���[.O�y���u��g��JbD���dCd����SB�((�|�ߙw��O�$��h�dC�`����^���=6�ԍTz|�.wV.ͨ��~�&%v����H�E���N�f��X�|�ڢ}�Ї��Au!�h��hU�ِ��j�"ҷQls�붼��l�ɖ�E��>��!z������)N)Ѽ'�X?�߀_��@4춍GԔ�lնq�iw��{o�Fv�O/����WZ�O���'M��
��{�^�d̓���׸V��Mn�&�O�;!�Ou�u�����p��*hۈc	^w{��Np&��#P8j� m���j����B�R��=H*�Zg�v�K{e˱���_/���~v��%V�NW,풰�(\�l��p�F@H�0�a�ٴ,���ʢܣ5�h���Oa�X$��V⧵>IO�����~3,�TR��
	�ч�=�
M֍�-NL^�ﮠQ�H��V����h�Ȭ�_AH��ҧ[��'�=�`��� ��meV�����3�a��:+>$f�XN�9g���*)��x�.[V3���-s�2��.os@�	�2ƺ��m����؂R����*_�~S�e"~�p��QgsJ<�}�5#�:�	����kL�k�>�'X�3�G�5�ǣ�nO�=�^O�D>�'s�Y�$"��*qȚ�i&���<�4́�~�[�/�$u�>�=��s���䰢ǟ-���]djB/�AX!\bc�&#��+"'��*��h@C����$eqh��XlxVHYEB    fa00    1500s�'H�26I ,u�d0�a�
V�U�*�c�\|��N�Ζ0 �y�Ǜ�2�A�J�悳��o��o�	і��w��7}��I����|��`f�\S&�eKM��xL�i"�b�?f<��Q-����Ð�BZ
ܕ�ܻ�"INT���0T�ӌ9�q�*����1~��1��6j?FnM��=�l��:X��c�2���Uz�\:����Y����C��Kq�G*~
��������B��_��%�"�i2u��M;�H�Yj�2����uб�^��ll$�@)��� �ǬDfr9�,�?�[����g�	\�L&��$�e�� ,�-�u��U�R͜��������;{�:r�8FL��*F|iN-��XX`��) �I�@%E�Fb�ֆ�!9��ݳ�I敁.hwI����z(�P�4�(�a'8+'JG���#�?n��;�$��L����#6�}m�r�X�_��_�u�Z0Z4:"}�9���l2%Z >�gQ5m��.k��J�=�٘�ѻ��w;B�r;K���~z>������	���~P4'M-0����w2�W3�=�牍��K(з�_Pyw��<��WN]nqC�ldd�vn�r����y��N�k�X�!�Dk!��d-S�����\��z���/��͎B^�Yd��r������Jmb�@��S�m�U�k@]�� �5��+S���)Q����:6�Y&����4f]W�֟MfF���Y2N�7o��pn'��)��_gI�&�>4�O��2\^��ݩ;чH����R��?kn�R[�ElbrR+�v`���n�(]�ϗ����-�^׉��a��]i��V�|���_F�E�*[�rk7؟�����
����Fs;��t"�Zx@8�Սr��x�j��?'�fQ�����GU�����e�3���LQ#��w1Z�Gx��۲c�Sp�WW�P��yҥ������Pov\F%�t]*lᒃ�A3�y/i��|���B֤����\���&4�;.r^q��U��������o��p=���On�*&z:�c��%����u��ʐ�:-�M�<�4�ʻ�&��)O,�|�T\��R^�r�E�vE�^�^ �]��%����ΎZk�$�O@�;��E1���ʧ�����������b���Ȏq�!�cQ�:|���"qt�Zm�`����r��8bv��W������C;�S��Iu�j�c<{�a��W��>xtg�����c�C"���6�[d���'�NK���",�m'r����6cFT��y�W�о�������Q@x�M�˼�}`,�Ѳ�˕��܏��l�*�)ZZ��ك�KF�8[ƾ��	�F��B^/ B+,'�1��>afӹ6����ea)L	����N�m9�m\�+1��>�y~���0!e}D+�R_������7FsE��\4��m�W[r;V4�����\�j�C�4��"���.�������cv�z��8DâAF�l�E�+�u�'��nhj���_���y-7�f}�w��dR���c�⚄w/�ͷx[�99'�'�<�X��m\����9a����!��9UE��8��J5������*z���R�"q�Ry�:�k��R���W���Fw�ˢY�'��G4�[���t��Q���b�`�Ye���ιt��.��s_|pmYL�h!/U �w��J#'�/J�s����"$l! �c6���e%��
$��[҂=z���LP,��|�l�p�H����b�SԬ��] X��~�2_ ���s$	Y�Wd5��y��&�Q(�t2pΘ'f��Pħ6�7�=�׉�?m!`�cB:��Ծ��pK����p�R4�ףl1fs"z`7�M����v��h���t�吜�5�q�Zض���,��8���>��.NԞ�]��Z������yO�9rq,����̾]�u:��L���
p�E9���sK���wD.,����|�4`:Z�+�IXd�XL1vD�90�W<`RQ���م��V�n���4)�ro�����w��D�D-"����1���n}�>��#?ĺx'&V%�e��y;Οesw!�.�r<��L��!��P�*��Ez��3��-�d,E�>�g�Bv��:Z �ob�7?��@djz�i$�G�R��D���8����K㢲���-�� %��� ��`L8�=|&���Yk)�C�rEH\ ����V�d7[�wxK�U:�*#�p��D2����iD�la��/���d��O�*e�W�g)��(M�ņw�U�W�R� �.S"�P�G���q-�F����$2lf��X��{�@Ɨ�D���ӝ_԰*B.�]������o[͠	���b�.qNM���.����U=�\/�����|o����fx�[֏H��\�7Kc:gq�l�^&���-��;���/��0�r����R�s�.�S�B�hF�R �cCWYn-��������������yQ#��b�H��ߏv�I�_,��
�n%��:v���`g�T{����M�������>�X���l��	��3�=j��>�
���Q�i�u��I�q����<�������q����S�Sӻ�L��ç�j*�ӂ���54E�0h`yn �B�{$���:цS�:��L��\�y�,��6elc�N���쒚�}.e���u3=�,��aLf�@x�MO0*)��뻍#��Y�9I(�����4�{�l�e�]t�t*9ˤ6;֞�g�&b�qy�G� T�����*IhB��8�D�����h׋&��6�V�8(A��v�?QF�v�C����+>�z.�|����<�k�:�3���Fāt+��������Ӹ��R&��G���'D�s�w��E[>�#m-Q�c�v�"�@#ʸ??��x⊏G��^��2ql�%�,�+*Y�%�ل����Q!|	j1�ڕy�p�N�U`��g&�uY.�Z.��w��Ȏ�I�@o���$+J�Í%�Ѕ�h�ߣ�<@�����M`�PĤuOb�-�sǰ��sB�
b@Ι?�� `7t�n%��)�ƍ"��R�#���a{�Z��z]�eW,������hg�2��2v�Eߕ7��a��}���i��-(�s�����ApzY8�.�p
�:�x�}��+�t�R;�U��,j���@��N3�^�똬U�%�u_]��fܴv���3�xK7��=�=<<��n8�h=X
��Q�혘�{�C�O!�1.�!^�dy�u����	�/ϯ^��=�3�l�ĥ��m;�'��96��e�2aL��0Bu�{�f���}�|��u�#B ;3j	 ���Yj��ھIɯ����7(8��Ǽ���e��Ye�����e
FK���)}:f������gcL�ܒ���E48l[q�龄�8b�фS���'TV�%_^L͓����u=�e��rZ��N�i��ϾbF-��h8����3qJbq[�Є x�������&UQ2u�ZhA9�	����`���=��gv����$<!+`j�#�̉�Ŗ|��D���h�Ec1���kdDe-�'��[�9�B�[��"Ȭ�i��?h��lȴB9v�2���$�/�*��@�8MM3/*����H��0��bVP�R�E��8���E#Ԩ���vv���!�L^�l��-��/�v�)iٙ���X������m�iTo�ɤ0� 	ȠkχQw7�0�73��x��]eT4u�N1�"6[�89E�Є}��Qv�?�����a>��y�A��@|�qar���%��4{���.%�X�/b�&P>�]&���z��6��'\�QtyM������evU���E�v!�dN1�ßo5Qc?L6&CY���cW��w��u�T��X�yۓ0�iP��|Sl��P����)�j6	XZ�L�&=td����/�4ߪ�.5ӉZj��Z��{�â���p�oH��ݴ���0�:���!S�uʷ�_�L�z�R���>b��jl{`,�	��8;V�@_y)��lv_2�!���o�>�*L%bw51�5�	�g�s~��OrǏ�)�GP�b x$��Ƚ���=�=�:g�����Dx�k��E�p_Z�:}����]�I�����7��F�뚥{k���ֽ�V�����d��Eh��-c*�o��:'شм���g��:��Kd���Zr�ܞqI��}IbԬ4a�{@3�*K
��p���z���8���^�ޥ�0z(_�*�ZUbՠ�܉6�8�x�������ێ��9I>��V<��9>�y��$2�υw㵈��э���W4�8IAզ�ıY�> R���-'�a�C�Vgrj�3�ӌ1��P�-�rtp��ɭsW9T�m �9���uM2_+�x4E1�m.5�է�ܭi95���|��� �/,��s����gfp�����f..,��&	�\����d�3t��.����U]tV�6f�b�wA�����ذ{|��(�x��:�߃_NCo���]sȾ5�?�SɏHNu�Z��1^�x�G�#��~�-­�K�4d�P��WO���~����=��Dr�}s��ј}�1J���CΦ�fk?0��K�Y�Aq2*�2��R���v�i��kV����E:�R����M�k1��;�����s*����,�nlJp��x#养⑴�됮�鯑�
�֬�t��+Z�l�tL��������@ʱV�}������a�auvq�)��boJ5,ǟ؀�yb��[�rY��o`2{� �u�Kl�y�L�SD��A��t$�:�.���<�ڜ��j�|Ȁ�1�/v=���"�4N��΅��m��@�B
�R|�/�(PB�phj�ڂF73���U����XO�M�&��.�s���0�E]S��	u���n�!�����V���Q����-{��ʕ[��[f�%�#߄�P�c�G���&|:�Rx�Ɣ>��������Il�<j�e���m���h����bg�W�4�8��r]J��tYt�hj��Sb��$�#�8�
1�A�\}����N�{|��-_�J���Ȭ&@N�3JOT�{�Lr�µZ�J���$��qiL|D��o�JpVl�u��8b�g�f����?Y{���Vu�g�P�&�;�t	?��1၀�������)E�M�A���y.����b�f-yW�=��Fʟ�[uW�7V��'`pV@��i���P|`�V{�U%��	~s�lc��������CWe��WC�r8xs'����/��I�z�@"�U�Y����YA2��{���gzv���8��Sh��c�٤��
�fE���XlxVHYEB    fa00    16c0L��ħ ���&�q���6��3���jCS�6G����L&Bo:<q
#F��w� ��w��"/��fM�u���g�.t�������hjr$���1�>�Lg���$��dH&O�*C���DK�58��UP�F>��Sz?�[!�� +�~�fͥ� Y����@�+�fK�՝f� �oΠ�,v�N����h���Sp{Qq�����;����d��*|�����I)z�>�O��7������;14K�A�̕H��9� J� LǪ�~�%	�eW�!*���㔭�@�И�5�����OlG��C��쪋ȸ9<<�t߽(�3!��}_IF��;r�0�آ�K[������vig('+�Y�v�������� {�Vmly�y�]�J�:E��`�
�����j�٘��|��kq^RK��k����w�#��<И-F���TEd%�8�����4�A�a��̫2���U�i�tx���(�=O���$1g�E:E�@�(~�3=��j�4:�TUiy�ˋ�0u\��i(�v�/��M�%��~�\ۭ翈�:�,�Xo��5��4�\B]���Eo+��؛�9��u�`<%�Y�N<Tl�r�*Bv����-�Yg�SYR���Ie��k�A�d�q�Q�/[�I(v���l�Kt�(��z�;Ν��|��@���<�K� ������aL��tQ؋EhUj��i�Gk��[?��l��'���+�\�	T='�1�������ܛ�	3��e~�L�]Iy�eH]4���Ȳx�ְȊ����(�N9*P�n}j���O�Cnt���o��y��ݿ�2�|\�ӹ�k����2����8�\�8�Ko=(F�A0%"�Xf��`�v��$�Y �<,n~�5q��'���4l3q8N����b+8Wi8�ƪ���l�YLO�fC�!Q�Ȋ���4�O������ ��X�?�=[7��{�W��E�G�P-ѱ@7�Lr1�Ax����͹Bs�*0�D� p\�*
�\9�9��Un⾏�<JR�'sR#K.��#4$�9t�tH�$w���>��t���\�b�#���q߆�/�n�U|Ԋl �h�7���\3���S�6�X�"@K��맴�b�m� e��4<�z.^=��G}�B��W�v�'e�Ϭ�	6��
��\W���X�x�b���9�'Qbs�%<��-ҡP�[����
!̧>V��ȁ9k�H�әHZy�A���J4�,p��仄jy&����
�q��70X!�"��>��eZπ^�o��
��x*��I�9��N��s�~�ݬ���;h�d[��* __������_r� y�p#��.Ya���Kt��aA�y�R�^�%^�LS����v��]:P��֐��#O��K�Ag�X����,�(�_�7Hc��{���p
�Ϭ[
�����&�k�6�T�����I*Ԏ�����dT�V��ʔcK�?����� F�/.7H�z�u������ct�m�$��u2�+{���v_dȷ.q�J�?�y�B�����L�E�b��T�r�"�E�������քM+�����&�P��sG�8�*�&��'gV��������m��.�۾�� �l�N��M��1�ëK�ҳ�+�4��
�tSA"��r�� ��V"`�5�����A�P�iϴBlFիK.0#j��l���`<��K��xIq�<tP�X"���C�)dݞj���F���P�'�'��Dٹ�͜ɤ4^h�����ƥv����- \i�#u��-���c@�Q�v���\*��ͽ�ظ��d]�*S�M��2L"��:�"�-��x'��7���ݥ�GK�v�A|.��I;� 	�E,0��ꪳz�dg�BZJ��s�N+^�@5ֺ�=�Z"��tL9��U�am+W瘵@�;�5=��LN����Ȇ�Io�P'��d�B��:W�-ڂ����q/1s8۵ڙ�����-�}��?1k	����{م�{�c ^�2�	�_��3oV!B�J�0��^J�{"�,s�F�#:<@y�.g� ��^S��
Q+P2�r���M�&θ$b���'��}ѩ1 �����!���z�62G�ϙ: ʰ�w��=l��{-�[�vW>O4�����ό�V_XԢ��,�'�ا�C��p7f��B13P8η.����u�%�Z�`�-N�
��q��ϼ8_����י��+���h\̺�L�s���D�1��tG>�M��OmD���r1�=�Ars�-�9���֥3���ԉ�C�*̻�_��������� �Gi�$��$�,��wa�<YRY�V�ۤ&��&O��kI�XH�u	�����6 �����頍��
�Na�ϽO ���gQ��]�N�v6C0��W�$$(?ky�����ѷB�xέ�k�a�����vOE�����%��A��MC9�^k�(]�.�A�[��o�0Ԧuz�k�UW��Y��#z�b�݂�t�	k_�;8 @�"hh�4n�냵!��qъ}�-_�ƳC}��
�uT\��s��Y�L��������7�DH�/CbM&�0�0����ӷ�%Y�'�ַ���Ce�NY�9ݜy���J�Ī�Ľ> 
g��)Ȩ������z�1���1����=�G�{��.�O# �b��=yq��@�
�CV`o��K")OA�䫅�Ǌ��ڨ�7Vt���(M�I����b�~���%1��<�=e��I�ꙓ����顖���ܞ%��?�m\:�;���j��ZH��KWa[��4���P����;r���j&#u�z��"���B.�h�h�`-�$W���V(J��*�J�'�w��MH�˂.�r:���!�S� ��	*���3�7� 0�)����	�\5���
=3]�����ڳ��PSh2�!���I@p�g���=��f��{����#X�h%�y\�w��h�u��G'äk�#r�r�cc_!:�N��NR<����H�=�$;��%�dxst�d��wm���}vhd@*�u5n��3&�A�3��T?�����{��t���D���1��抯�~��X�a�)�e牚����/��7�BrI�8��.�Nʆ��sV}�	��R���G`fv���-7��<��S{d"��~d���2ʈ�����$1wJ�(�0c�������/�X�� ֠V��Ğ�m�dYȒ��N����,�_���3#�ƪ���΀5�pe&��2�q�u�H�6��.��|�˓�?q�e��� ��u� ��N٥�����B������~��Fp*Ym/��E+j+�.�Y�q�Y�
ciK�q�^\�6׊������U[�I1h���'.	Đ�T엱N*�tA݃�LP
�p�R������D�+΁-b��&�,�<Ai<_����cr��X.�kZni�zk[�GxY%)Ừ/��,ޮ.�^үVX�E�c
e(��.��]!����hny�`��)��&0oR�~1�o�`��߫�H��j)�a��J��s��lH�4�c��"z�z{ۤjB�y��y2��T�Pg��UL��m/����0�G�\�켓��ҿ1���<.Pr1K�t��	�Nh�AJwcc6hM��:�Z��Dp\COh	���/�O�%�>�ͺx�v�VO�"��2�^����+^2������ٹ�^�nF��M�{��|Tɰ�� =���7Ʒ�K�J�ޤ#)g$�O�켶�*��$_���
��sA�ٔ�{��Q��Ki�Oh�g�5�K��oj<��I�<A�1o��z�GˠQ�+���b�=M�E"���f?r0h�=`���0����_G�>�Ǧ���iE3c�hҸ �,��`���H��v�D���6B-��3��KK�=��Z�V3Qr��Y����Ō���1:'R`	�R:k������6Ǚ�"��V­�vl�2�h7@
�R,�0p�l��#X�X�+���)�e贌�*dI��y��Jp�{��I3	���oOj]^pU��Ԫ{��΍Ov�VM����mo�Ia�A�F�������Ź#��	)=w�^��<ȳ����8�2��׳1�[�ա3LY,"�=�KKU��"Kɏ���1�1&�$%��������k\���tJ�F&�o�~�W�Ėc�j}�^6�#��)m�"=\�fj�/J��9�C�`�1u#����֯��q�����t�+�/6 ��ޥ����&ra�ѹpbOzN���t�O Man��b�b*�=-����K� � ;8��մ� s��n+ �Y黰����c{-���<c.�r\V^��=�s���x�Ǵ�&r��[l*�gOL�B�فGI��΍�9�$Ks��)ɖ%-�� B�:!y�]��
h���_.��P��aZN����5u	�]���0�j�mK�'��.�+5�9��Y4�1�07s���n�E�zb���^��:6�s$L6���c=�E��C��L;5%[�.��&+���2 ��#o�t�����s'�� @��Ǎ=�����7�1a���7%lL�eu�n\Y���9ڞS`��o�$��솜�w��i�}G�P:���.��*Nu��8�������u�Y�M�ZCYf���� ���jO�mQ�����tZ%�	��e�\��{-����M�b(D����0������B9�Ɍ�Bl��[���z p~�({8��z�P�rT������
�넝�� ��b�z|�uѺ�F���v���WlSe�u��>�V���A�������C˷���g>��+�̈́�ⱺ|e���)���K�^lΪ�9�V>Mr��i�u�� .�C�ܞ�����s���r��Yݼ(�9�ŷ��+�-�]��Ys$o8�8'�^���r�ݺվ�I���9_+����J@��"�D���Ĭ`�'�8�|��τ8�� �d���]sJ�I�jkZTŦ��B<P�p
����\���eCH,n#� ��3��䤃��&� .�qu���v4�=8�	�lK��/>����o
�>����k��F��Yd��@x9V|*�G��?n5�+o�̈wޗ�����$�!�̀�K]���������Cv�#~�̅J�����(qi=e/�M%���3M��9�#fD���Z����8]\)n�H�-�f�Y�pJ�$�`F����Q��<LʧӊC��8���멋	(���h���i>�U�`����E�5�HdǞ*s�ϭJ֥�2�ѥɠ�
7�̲#t�iW���J�<u��8}!�i#0B���s�]R��~�,����+�Gݓ����IBpM63��H�ì�b�&�(�ȷ�m5geDu��K~�'�S|j5�nk��6 �xTCM��㉟����#�4�	���3�{܁ M��|�A"�#�=����Z����#�X�[���SX7s(c��DR{mw÷���/JTXh�/~�n��(����-���¢����ii�E}�t��/W��ﺪ81'�p�WR?�{l	�&���Ϸ?��r�݊=	/�e���AR��{~��V�<U��֖2zj�z��/��|����e�Q=���?���{Y<��~�+� m�fs��$vE� 1N_}G#��������}to�vդ]Р~�K.H������c����Lh�8Ē����R��WȨ��5?4T�&�"{��F�Z��Y�)+*��-�^��E�:D[�'hB�T������8���stnW��ꍶ�F�s Yr`f	(HҐ�%i ⍱u	��&a�Q�� ��.�֎@�2g�M$�h怱XlxVHYEB    fa00    1740�H�@u���q$-�#3�K��p��S��+�I� 
E:�&l܁lc��22��%����L4�M�͕ae�doq��w����n���GƸ�F�u\I�V��%�;D\������4T���n�\L3@0�bdb1T����n��^CsF��O�qCx�f�	��>��p�5B&�^Ac%װ<A?���&[0��~�>L|Wx�8��W}st�s����1�l�n�*�GQ��0t;��x�����b��yx�Q.�7�ϛ�"�[����*ӯڑ����N2^���(M�(֤?x�(�7��=��aP&z�hu��h7��s�䖸��D������������x�>������?U��sphް�o�>~D�B9��`�Wd�V���#�^��Z�i��!�*#`��F���L�Լ"�!��23�
�C0 R��u)9�|%	�Ԍ
�w���ki: �SR�����C��fI�bw����T���~Vt�m�EI�KY�/��Y�����t������Ws�1WȡfG� ay�O h!��&�a�8;[r���?{)>L3u�a;"Wfפ{M!��8\Q�+sz�;G��o����6��Ԥΰ�ʔ#�#���QWڟ��Gw�����W�b���-q�G�V���~p��!)�1V�W�##�8���Kt��`Ԧ�����M���{imu�Gz�7��a�0�b�s��?�qg���vv�X(n�rƶfO��njL+d���T��A3�6L5"�']D	���0퍝��V����G{m=����bbX��
�\�, �a^�����B�{IX<m����1G��t�r��_x�ҍ�[7^��Z�w�B;Q�bZ�n�g��3)�>Z���+ׁ������ӃJ�!@ ��C������yMP���]D�f��1�J�fd�Ćws�蝡J4\�!�fQn|�Z���:��!�&�($�v"�JΒ�%_��}4�/5�4�zv���G��{㏑R�~�{K��2���E"w�� ��a��{����By�Q��a�"�^qI�7� �0��3��np�״D�v��r�n�o4�w��m�c㘮8��O������^o.�\|	�w���$,��N}�(=%��}bXasmW4	٣���rZ�����o�+��)�b2���s9X����I񅷁�{��z'(�oOb��3��R�Ӏ�U�4�%����:K>Ud�~�(���6k�~
��\��T�Hi�����;�����\��C���?Fb�Cg&�b�Y�f$����/ ���\���a�E��*��h.#�w��� *���w��)^��x�9,H0$KXQ5�<f}��_�>б`(��J����q+_ɝ����H�tE{��'�?���Z	鴑U�+�l�x䧄��Āڵ���@�je�W A0�s$�s��Q�%��l�L��$U�.x��_�	�!���� ��A��>�Ғ�;b87����=p�{�ΤW����<:.׵��͏���`;���&N�zl�*��ؓ�
�;��.;��Q�#��ֱ��ß
4���r�:	YY ̯�#2F����Ԃ���`ס�KWV�ư��j������p��.y�n�%ڱ�1\�}{Pژ���#�$�[���1�*Z�{CB
aI�b��o�G��*��A	��a���CsH?B���3>�ж���
S���;��j~�&p|O��}3�/N��:�� @���]������C�qx�i�zE�~��&Ni��R�\�s䱌�E0�萣m�}aw1V�j�� '8t�E���NMZmo���Y���e���"���S_�f��=q}� �A�~%�/�V��"[%�|\��J.ˆ!A7hPL���e�3�-�1��J��(�F�UH��Z̎��=�U����my�����<�5��XD�/��BXɣ�,�����������O7("�(nZ�7kX��LS#xT��
��b^(tO�l� �^[�2�n�ߜ�0�u[����su����qnΪ��F*��;Y���K��t�f��������Ix��NS�AѥGS�	Vѧ�}+uB݃n������L�ݐ�+�"4d *�$Sr���C�0�eH��K>q�I�o*�7���V
eWƬ��H��i��+a�b�(�ŴM����XH�Ĵb�a��`Ϋh��Z�E8�$�&I�hXڂ����EWk�$Ü�Iz�E�\�o�=��������h���y-p��K�٦1�g�b�M(%sfz�E�7��tM�0E<D�?�>C�%i}(ķrٹW��4?a�3���p�7���n"�b������})�KK����n�_G��Y�A���#�� r��Bhu-U��3:�ՄY� �g�3e�#���xb�F<� �6��-*�^bPl�m4�O�q�&w�����gc��k�I�[T�pM������w�~�B�Dk�	���ř�so7����q�s�W<'�+��	�2�8��>�F2��_��>L=W>1�D�/�Ar���޴�ȫ#Ew���xFh�wc���V'��n?>e�ME
@7̩i���m/:4tϚXZ�?AAx81���\��K	��In�DLw'O+|
����LQ�7MT�椈g U�U�6-��q�v��wԂ��Y����`�*����ߕ��ȑ���ok�q Fߏ(��jCD�^�oB��y�=�;G��#xgsdkK/�>�J07B�������`����M:�]*�Sٯ\@��64� �挌8�@`/p�^z2�x�������zz��;�M��8{u�]a�`�ɒ&��&Շ����f����)G�����a�߷�M����:�wNc�ʪ�\MEV��x$g��l�.��Tr����Dޚ���t	Q�N+Z*���7��*�	x��o�%�� ���t0���߂���|O�( ���WQ2�u��Z�NY�_��:2��Q��뀺)B�54w��HY�f���뵸��<�Xw�ͥD���o�)yw�>ŷn�������?��5;*���o��؛{�J�q��3�k�@b���}�
n�R�vXV�1�I�[�ǬJ@�����5���-����aMih�:f�����~��t�!է���5�����_-�����8E��|c���o�9�iNS'�H�\^l?���i=YD%K�N�k��F�\ɁR�5_��]��YO�hߔEAܻ� �����|�W�C�|O��LIb[*Ʃ&vw4M��!:��⁸���X���������n�=�pug`�����Ƨ,l*�@8�D��]����M�PH�v{�,��M�"��v�r��W=�'��fsū�u�����¿�"�*χ��x.+*������k=�� ����6�{�!0��x|�w�f�>�~&����Y���&)�:����;I�S�Ǆ��]^Ka�{�" ���n�F���^�Ϩ�_�3�q�%�c��&���}�X �9/bc��+���_XC�u�gC��(����$RE28\���#��;R4���ىIӋGs�F���Z
��X �7٥ߒ��|{��!��yҖN$��Q�d�?f�b7��!���s	�{&���҄$�A8��|�;c��ͨ��� 1io��ak�J,Z�+-���[�����&&0����.c��݉��Ď9��`�
���v���L\w�L�u��8���R��wi�h�$�����t+�s�0Ӻ�REQz�~��(�[�m��\G�W�pk?WImb��@|:�#1_\�U�@M�t,���zG0�@�ү���	NYu�?�IG��xh��s���n�M�)H<Mn�Z0�>ҕ=�b\ib87�	��v���wۦ��`����,�f�z����J:m-;�/]��
��2��"�{h�Y��=����н�v��/�v�c�y���N;�����'�u����䱊��=�:��e��gښ�P�ԑ����	�=3�Є�c9�>���4�F1����z\C��m1;��Dq1��oL� �jM-�@S�T�Xf�Z���nI�l���{�,�Ӏ�6�9�t���͏�{�Fݻ&%Ը�c<tk�V��'��~����X���N�p���ON�4��O��2_�"7�G�>������"Q�@
�i8��E�x����'���-���♨�������e��@�{E"R�r�Ivc=�*s �4K�v�2t3bT�QB�F��$i	�g�E�L=���v�O�:HR|�=�4u�YI�nR��^(�^n������
i���_E�tb�>Ԍ
�۽@�]׵�_���)�>��*���-�h�1?��V�o���z��;r��Wh|�U�l>X'D�EZ���K~~�`P"�c�(�d��%t��e��$�����j�'(��S-`����3 T���W�o!G�b�ĵ*���T4�A_�X����r_K����Q�+@68��q_�]@N/I˘��_(���m�%'ZU��	���f�d_ "�` ��b�]��ٲ�ͤN:S�&(D�v��EL]S���G	t�1�?�T$����� �IF~��%��pY��7�![s��)�F߼/z��8����' �6P.�����������':��,�t�6�Y��'�W 9]��aE#�\#,"��;D�R�Zǯ F�����T`i���9��:0ߺ�&��H�%;��_U\�o1@�2{�S�*=3ck��Y*�U_PJ�����a���˗�{I
0]�qAr�e�ҩz���*[���V�\�:,P!$t(k�eF�`u��9����0
j����
�Q�%�w_uy(��$#(K����<�e�At^KVL�����N�W��F=�3w����(;�-k���	�MH���aȳ��9��`(,W]Ď����ӾۑW-�oʿpyT���<	�G���Z��ي<ȉo�7�?o����a7�9���K�ʁ�/�G�������YD�n�0=���n)�1�RO��l`����	���*�zڮ��<��-�cX��R����hJ�(���>�@P��}P�U�	�}�F�>����{�q�{Z��
�K��o��S5U�N☶���2�a�-�	���X���Q}L�T)QL<ʷ����a�8��+N����M7DKcr��t��2��i+¹��������/	$�a�M�� ��i�j��{H��v��>;�E��ǃϱP��#�?[J�������Fw��G.�H��V�ǧWf���0� ��oľg��{��������=�9&�"�L�/H���űd\�������re�[��^����x��_���R[Wp���K�~T�u�uI�DD��0��Ҧ&���p71h�=?2$���L�8<X�^E���M�iM=`|�A_�|�R�'p��^�-���S���{S⪘� �,�qWӠ�W�i�zXg����~K��w2�^�04�����?���R�^W�k�sh�<�l�?Lq��&Ą����6���� ��ƌ�'����~�Q��T?ؒie��m��D��(�&Ś��&�����'C��`*���%�\�W��"��f)2F�����	紨c���m,oT�_�E�����!}2G��0�2��̋���*C�p憎F@m���1���Kv��������M`6��x���b^Me1aǕ� ᾕ҂A�=IaEhd�ݥ^%H)���2��9�����e�C[�/P��s�u<RXZQ�;���9����!
�&��#܈͹>P}=�w���=XA0���>�BqI���Z���4I����+$�#�Zw��V���4"���(����kUv�Ō�|e�Ī{����[;�L��݁"�,�9hE�+Su� �)�j�Àqx��[��nq���V{������l�i�"J��>X�ƥ�\�/A�}�%J��4�#j�5���XlxVHYEB    bf14     c60�)�#e�Z�'��_���Ag�)�8#T�#�����^�~;��v�eC!Οs�DK%Uآ��`�T�{� 7�~������A�^�f���)��T�՜�Z�������;��TxG �6�m�4�D�S4ni��i6^��|�!�t)�2R��������X>�~�����	m&O�XO�d����z]B�c�&kӾ�^�ĐG�|�$=*Uy�����BD����}�W���+^�g�̉� `����y��|R��eV���tc~f)��v,��g0�
��r��wÆo�_t˪Ƀ��Q�v������Xڣkh�qҊ�g�C�)8$/g�Pyoo��鋚��p�:U�~���H���8���p�
����d�[�j��	�W{��P��!g�����"���`ҫ�v�vA~C�C�X٩����GygHsǚR������w�l%-��!={on$��J%��:���5;`��_�"�X�r�b�
�s��]��}&@�VU��t@́�|�J���G�}�u)��e��jݙ�[T��>����s��	: ����E@w �`��W�F�@}���0)n(#�.Q�	t`| �& �1�9\�2c����� ��z�#���dXÑO}�[Ë�oM(�5��޽+[�V�y�[�-!n�Xd��mU�W~� _� �R(�_����ǡm�*-A� ��2H`^� �·Pc�_�y�ճe0sBZ��Rm��-"z�y�!ӭ�����@�IZ!��t���4�a7��J����/Lwۂ����xf�ɮ*���PI!��Cyq]O<�W�o�����!^
�E��P ;䬙Sc9Xs����d�� �@�m�rS(�L�w�eF,�)����u�ȅ�l���f��P�0dq!��*÷:���cp
!@�y�CT��
��,�;ѩ���A5A~�2��K.��S	�	%8�/������A��/�E����4��R+B�0��(���3(���`v:f��"�]�^���Q�Z�9��:�1�0<���Ӑ\���u��.t�|_�������=\�H�ʅ�~M
`ߔ>�T�6�|eW<D}�*��w<8�0ba�k}'�U�����s�2���cZ�ii�2k�=TH��Q\�L�]�*?�֑�xSu�
U�j���8��b\��lz2u�xE��&f��&X�uIb\�G�B���ѝ� }�P��7�*�̻���ؙ]I�lq�������OS�=̏ȽXN]�� v��M��ps���o�1��Tg����<[�H_�g�u��Їq�?Uz�<p+Ӑ�BBI���NWK/ϔ�����g�Y���h\��W�aO���
�ba��!�|ᴶUz�>��#��_���z���F��y셏`߰M��E�m�
��A��S=�0)����}�yr��C���t�4U�{��y�����X�m xX�I�9(�:m�pk��$��?�>���a&�6�$Ki�Y�o�_x�ƒ�rj��+���b�"ZP�� ����-Y��橀u\�w�d�r1���6o�p��%��4�]�`0>�fR�V&*���K���\,9
z21���E�3��l}�+4�#��#�Ԟ�ۍ�=�1m�$� �F>���<1-�W��m�0�B�A�.L��Z%� q�?ٍh����gl$���t���9��R[��؝@F�1�2��ݑ��� ���޾��nK��Ɩw����������w2�
��mIyC���S��U��]�×�أ �ċ��P�9��@��	<��4Y=SLl/��l�?�wE|��>-y�x���B�uԽD,n��\��9 s.	�Q(_r>��XG�f��Կ�f��q��s̰-ǖ�0�{��}�6'�
N�7��rC��)\%���G��[Aޓ�(�)����g�Z1K6yFE��MĭYD����ϙ�
U����r�-�ݗ��%&_~�p[h^͚�E����nD���s����^�!��3@g@�0���� ����M�����;=��r��@.ic>��F��z(j<�
�R���}����D�d�{$�R����[)NK>F��^��Y�cI��c	���ߎ�-N��
o�ڌ�|��~�Evoc�Zf�-��?�ɒA6�Y��4:�<�S�:��[ͩ|ݲǴ�,��O�\Î���3y��Є5e�e";��;��CWXw����n�˶��[x�#�0q���6�2#6�z�����P� @X�c�&M�ҾO�b�~�=1ݧwd>�h�l4%�^�E����{�&��qcs�r���?��1��5H:��ow��[~�G�`����ϰ���l�O�X~� c����Ҵ(x�:�Iy����sP��O�o�b�O��Ѹ孂o��R��q��.'GO۾�@F#��*߳k� �fjFY�uy ���;����8���<���8�
���"UMU�����"��6K)�d��4�K�8�r4{�R����.��\�j 㧇^��R��U+����ɛ��-�=-�����;obΈcm���#��:C��*�;���3�!�����l��btuξ\��7��������odq�������y���J@i��ȭ�=�n��RK��5���"�A=����Nk��~��o+�B�V���uY����X��\������_�j �9��Sp�7���6k��M,u����ظ(Ԍ}�����L�s4���[��PU��[d��o ��#���4�vK8c$`�����:`WVL�ב��tɍ̆��(	ul;慛��r��Cԣf�g���t��y��]_惻��&S���W�sӫ�k��`�����G����i�$v!��
�0�g�#$kR�#�'�T�Th�,�|-�U+v�)u�:�#:O���9�������#SY�UY^Ԏ�t�O���_7Y�׃�4,��'N��ʁ�Q7���1�K��Tr](�2�� �ե��A\E9�<�]�9X�u�}-O�u;\3�����g�y��}��sD��#Tg�6uEvqa[��������d���-v/&�F�F?q<�A�̒�r�Ǆ���U����4��Bu2�A��q/��]$����3 �v�
Y�x�)�c;ꠅ)uT)��]����&��7Etߍ�