XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���lªB�q�`�e&Gl-���8�y���[��籺_5g����Iy����S��1��Ț0�{���=t�ƖK��U�����%��w��^0�ώ�H6�������A�:Ի��Ļ�z1�u�s��J����^�[��u0T�la>|�c�1A�M�;��:Glf�|�p�润��W��L������Cn�w黦b��A+)� �B��c#�'�Qk�]uc�yz�)d%0�?Ӱ�7����5���7qϾpD��+�VW��j�A���)@5�����������m1�<���U�T��FJ  �-0L�~=�?�W!�Сۑ��Z��0=;����;7��E��*���x�p<+TKv��,/�(��Hu�su�j�����u�.��*U���Z�=<�	�Z��a:O����NY�]���Lt�{�r_ ���bډ�o{/���{$��k��lw)��Jh����,h%�`_+gt�.�b[�����U?4��	`إ@�U����u_��C09���AS�Ōb��گ���2��o��xH�����	�$� ���˙.dw�j�u�)� :�t��2��e}���_� ���PoX��x�g�m@q�V*gy怉���%R�-�ymCoy�:���|"�ԏ1��M��"YédiP�峠�$�39�����wd+�7���ېSd�q��2�3�� ��+�h�EfRS4��l�ia�I�&%���B�Kp�U�=���Pˢ �(�5�*^�-�5<��|�XlxVHYEB    fa00    2d60��R��������=-	�S��®fMLDʑ�!>�0�l������G(��+�1ی���h�4�@_���H�<
�x:U	/��S�(uή�\M��Ll�/�D��߬&�ͷ�M����I�*9�96�5#��
ȹ�-
s������h�Ζ������R�&#�S̼gc���T�r�KQ�1/�y.tBW���Tf����b~o�)7)X�R�Y#rz�E�7Qe`Tx#X��Sk$�'6��(��J�	c�ү�.7���k&�BmU�;����N���)���M��v�����ű�Cr�G&��+����*�@Bw;�C+=�jSzo[��5�[��8	2�8��C���k^L�YG��{��P	�ǹ�7bR~�]:�bX���Y�DX�"]A��.}|!G:�� 2a��o�V{��盵����Y�U�8��������`FŜ�[?��2@�dB�B�� ��H�j�#���]�5Z����P`�&ӕ~n�fY�@��������)�۾�|�2��
I~��Ϯ@'=(OF�n��ͱYk<q��`6����a��c���2��U����p�
�[ކ��hX?�5.�J��!0;�Pu��[2`Ԉ��c��5�#�Ϻ^��9������N�o��i��L�W��'�|�v��8�/�c{߉R��ڿ���7r���B�X���O���6���>����_�X���!^v�O@#����<j����Ka$~y��(~�����ÊTƦ
V��2����~�X�i��E�: ��{],��OI˼�7���˻�V���a��/n$�?�G|ը�V�,�ه�FS�
�2�	�t�LO#��h|��ća�.G/�y�Vyr�k��qx�5�����~?�}�rC��X����:ɸ�!I�2QPԀ��}�(#�Zd>��i�9���1~o�mA#{>������?���Pk9�z-v3H��~2��z�y�R�c�AҒ���-�Y�FP�3 gJ�L����_�D�6'���{����F�Ϻnr�(/Q�m�{/����勁2_'��9O)�z�����8������p���vH�cQ1P'�YҖb>��y�8��p[�� ��:c����9w�a�.B�\B�*;(3��ie �3#,���r�8"~F̅��  (k��u`2�b��.\RW���Ɛ<ݑ�g��ZI�a��2~�}1�j�1�>�UV�6;���t���Ǽ4��"�H�����D�ʺ�ȷ�7hي���03�WN�1��C�P,7_0�/Ŵ��q'j��жx��y��}o���{!�
u�T���9�xxy�D���H����~��[�NE�l���W��4%�":���5����m`~��^?�09�5�ٗ4A�d�c��W�.�L�#g'ux��M��m�-tרּ`�KS��ܗ�0>�n�e�ą�^ju��@X2p� ډ�F�����'��;�z��EtU�?�vS�o=��MZ�"A� �Q�/���Y�R���Ǎj��⩐iQB����)@����p��̔�D�_�t�a{.�V��.�S4Q$e[L6�2f{ˈ��5e�+tII�d��;tAh'ťcEڿQ�����;bi|�e�7lv�_�?K��%�����T�ڕ�YLX��"#�=�.;0Ɖ�U5s��w,*�5Mf{w��TXG������@Q!a��_7�g{����l
H`j�;�s=�O0S���p����_� N�d{�"�]�U�+�7��a*��]ZT1����Yr�����'�:���kD�)��d�>�T	#Љ���ZXV��)5(��(�'���4tD���ѿ3�u�[>	��<��"o})���xڿ��ji����~�{�Mh�b��x.g��JO�R;�������D#���n6C��o�M��;�h���,/�L�<�f�vm/0>�l�ŅS}��)埝瓕��K�<�rGVu��!���By�:�ֺa(F��M����C�b��jd�ɪ3
'����߁73w��������SnF 4����bf?|"�lGŻ����i�7t��2�W�k�A���g��?�ߝ=ۑ|�`�Yv� }8�?�]*C�h���U���e:#>�|(~�0D~ȵL'�r�sC�U9�3Q�s���;���*�����Y�v�<��͍o�/�� ����0f��.�z��sƯ$Wu����t��tL�H��fؙP��c�2犢��,�כ��'�^l\T�l~���Z\�����6��QG�W?��ڽV�p��9����+Bu�;�E�''�#xFrv�ė�w�e鳋��n�.�e'o�OHx�A��i�\\��}f
�2^ң�Y��5��W��)G儔K1���=A?���4��g1����;��H*�����S��ڍP�;;�++����W�dS��<�%Y��3w���+
;��d��Ãx�'���s�:���X27K�W4>���<��m��_�{ɥ���־-��X���P�7�?M�����T����	*\���Xh��]b�4�͖���F�F��v�q�]�Id�`�N1��[�P�3i���ii�r�؏D0SM����W�U�����M���Ħ\�>5U�Pzj~i��ٷdH�(���#�HYH�u�%~��th��T��f��A�>.B)4d2� ��x.��8"�>(���W��-�g�S4��5�WϞ7��e��򋮕bRP���Uq����k�o��:rq8$~��*�-��f��q�ҏ���锪��?7Zm���ڶ'��
�d�
��7���y�=�3��\a
gd"� ��r��2�b
��K7
�0T8ob9�B��#(`�'d�Ⱦ!���a�^����}���L���?��E�&��c�$�4�O��aB���p4�ߟ4���"K�w� �ı~\�>��Թ�4�����׌�T�S,�Jo�zH�ڭ���&���ut��K9*(JU	7;S0�����0c�f[���+��T����[�|��]�7�C)�==�0A�\�S��d4mT��ʕB���,�A[F�1�;�E˵	-�i+�W*��"��2�t��.X�%{�©52.A�Lm�z���<���?w�`!��%i�;�i'I�t0J
Rʇ���|��5�X����fY*I��a�Ƽi1Z)�����MaX�Bv`�n/�yJHP�Q�(�B��Gl���! D�����>��7&H���"ܻ^:���A&v��9s��R�e�ɨ_��W� S�I�����]�)�� >s�c�>�@�o��9A�S�E�C�\�C�J�M"A�����O5���]!n/�A_d	mwy_�+� 7�rZ������Mf$�*_2����35*���8J�Y���_$\��3�[D��%�D���Tq�kC-��>�Ŏ���"��n�\Ao'���"e���N�(~>�Y��wi��a�v�'��<�{�l�p���"aV�~Ѭ�6�5Tb�)��W~N���!:^:���_�	��[�C�?�ό���〸 �K�d�Ė�����:B3�)Ӭ%C
���`V�W�z��������8��E�a��D��a���;��T��^����݊/;�lX�����ꕐ��Jf�=3]��[��,W�w�X���N} �\7��N�x�N<����T��0E(�,����c�W�����7}+��������_ޒ�&�Oz�i�>ܘ�`�6�%��]���:3��!�C�q�wb]C�IT��lZ\Cv�j|��{�	q�<ϾJ��9�(�Z�J|(3�6-�.��u����
¡�T`�/s'x?�-<�^!�>	x��S ��Ժ��r���X!�2��u<)`c������;o�H�B��%$'���=;�?���w_)v�kJu��n�(	��O����/|�f�R���u͝�]��?�[��n�n�{q�8�>��~M�ܩ9ǰ"��c`���G�X�ɻ˜�ۡ������۷Z��I!����N�U�<g�4_���)Sd�h�?���*@q���u��&H7�9`�y��w��M@�x���n��"��U;oF$�WS`O�d����U��]�2��x��are�3��@�F���%��?���E�z�?+�;�����v�g�Ƽ���XV�-k�+�e�k��`V��0 X%�n�&���GBއ�ݜPo'��)1,�-�!j���M�Ճl91jP�GƋgW`#���6�R�遂A�6�l�#��sR��еdt��3��b%{݀x��S �/���,VJ��*�)���8����RE�KZ95b�<h��	�,��!�;	���D=u�3��&�b)d��^9��HJQ��"�AǦ����?����	�J�i���}T��� @{��\ᄌ�5I��@����S}�2%Y��O��z�t5���a����g�Q#��m#A�2~$�ܳ����	����>�z��`,y�l�pOǱ��6	J?`zc�'�E�:�m��sv�vl��c�+�q])
���Xj���C�|,T�xg-�5}�4�K������gnl#O3�9�c�/��"���]c�M�X�12���Oe��+[���<b�x����:����4����eǈ��}#���(&5�4��wj�iMc�>.�����������p����)��'�L-�Sse���ƭI�a��d;�T��Ǝ6o�.�� ��!�X��M�Z���j*���{�^�XYB��S+�F]�Cb�$Z#R)��I��e1Oc���9�)��g<&!.���gU�^W᪤��!rj��sĥ��gn�2��Q�g�"jie<�s �;1q�q
�b�f#���Cg����Y��I����W�g	x���1�Q2�y+TS���ޕW�u�c�dQ ��T�eH�=��e�u���/ 
-��:�Mﺖ7�_:Y
֝�ig���l�_�Pl���j�ף��ቲZ�0:���f4)��F�u2u\����q��fH`u*�#_���z���\*���v�x�5�^|�fŏO�Mv^�N� ��^�7�9۲&ʔ*&��*w��_����Co�{J�b$��A#���I&�d+礝 �Y.��S;^��h)�.����L�v_�ۿ�Zg��6P��ٷU��ugѦ�B������|�qb�����&�����-��qm'�I6>%�v2=-���=�۵�l��q�g��Hl����@�`�^��f�4�x�� W�d�5mS^�<���v9�0~%��}�*{�;*j�Dp7'���Z�hvC)Y��b����X�߶�O���i�Wk1�ϻ�m�Vi0o"̛XVc&�m�� �Zj/�n�j]�&C�_�}��D�fNU���j#���S0�G���ȷ�̒@fY���EUj��Tr�T�Q�]���[������p�(��+Q汧�j|mYA�\��d���ŀ�8�E�:��U�+���ަ��$���A���;UiBN�9��$�)w6(<ċ2�Y��m�֢c��1>&�D�㭖�Jс���|���Rh�v?��T�"*�氪>��2�	���_�g����9?�`��3�؇}c��֥��>��L�m�h�6��1G�c~΁צ����'/f� G�p<�2�/<�!�)R�*�X�C)p�zI�����Ĺ�ZQ�/�p���\&�����>�A#v%�*j���o^}���w1��� u�[���6 D���/H
V�F�S�h��vQY�]v
*�JŃ�E7�6��D��ƪ�À�����p�<�g��Q��c$��MY�7�����m��4ΒB�&�����M���v�p�����8_��8�A�pl��K@��[����L��`�Z���磐�0����F�+��ɺ*����zv�6�cO�����Z�i�����[�������7`7
h�Bs/���<�B�v�p���#�C���{����$��&�K�4+\<�-��t��Wn~��5W���A�~��6����[�����J�əbN�[S����UÚ0B�`�x� =F��i����JK-;8:���v�$K!��+%�eԭ
%L��c�2�Ӭ{D�� 5ް]�5ل�n���.���ŗ��D݆@@"C6x�t��d�KI8��`Z�1Y�[ϨhKt��s���,.��ʂ��	4�h�vYTs#|� �;[|󏳖&�8�vyj�Ҹ�ZJ���h֟�Q=h of<,�"2@c��Sn���)�v�g�j7�����UL��+�Y#Wq�r�n�S�{Lu�M5���f�f��=��@
n��F��q���2���A#�� "9�ˏa�u�I±�z��8��Х�ca�+�>:���	|Q�Z��-(J�Q���;w�B��M�W���3}�S1�KtcQ��=\��?��+�Z��~��މ�e�|n��h�{��a*�c�%�nlČwג��@��|b!���lU��U��R��A-魉�i�J�dp@�;�n��p@pJLL�CF*r;�ڤ�&\�&M�c��MU<W�Z&'����-u{��}���%/�ot��D@�+�H�r^$����Ll �?+5F���:Y7@�%�X��-	��^���T�Q��0��nW��[�sE|����-"�F��Oc���ŏ��cGXɿ�iÆu/�q��k�k�¾a�$2n>��oe`���;�[���guE(��� ���D���$Cq v͢@�?�IS��oP��A�9.*�Ԥ����V �J����)4��k�*���D�%տsa�ç�f���\� <��}>6�m7TPvq�'+��
,����8�=_m��-|�!�,F���,���AH�_OkcJ���YW<y�Vh�#t�ǭ,Q��Fv�ï`���#U����5��L/�������Cώ��|V-�O $�����\m[7gŹZr4ZHa!Tw? O�9g��l���y��lvݐ��U]t�����y�~�8e���Qә%�h$�� 0U��}4g!	�.��rJ��L�a�$j`����$�$�����>j���'�crN�ɥ�VZ$���gBS�]s�a��3*�W�B[��g�\[����ѱ���딥�B�Z/)�����qʁ7�yvn�Qv�DN�a���m4
�p�T폰�Q��g��`p�	iA� �#���{�
���=��`���8�����)q�e�匔�sX)�=@�~���ٶ}ځ"~����.���̕toA�X��a��А�u�qB�����H+��+�߫���<u!��DИ��sT�o��R��L��w�հ4��$g��m�5���N�{��B���D<[-��xBL����c�D��10;l/wr.�Wd�9�h�8:���ƍ!><�8��"�Kv���d��碘�2��R �yy/dN��~�dp����-
���TX�A��mW�^�%k�b��g��Fݖ:��ݯ�
t�T�+��/E���A�1eV ��(�[0v�R+k��Z��^��{�a���|[��l�N<���#<O�W�50�� m��G1��:�ý�E�r?ՠ��*d���a���)��n��E�Q�K����G���)�#���ד�b�?�EC1���vȃ"4D�(�0�e��r�V�,�-��*��hǮ�� X�&la��;,�$$�1,?O�"f	���D��S{��$��w!���8A��6�����/����:5��c��0s�����ta�2�4�l��a_D��i�0*n��U�9� ��|�_�Oݴ�H�{�.�� 
B���~(����4�6�sn�,ܵ�����+,!�q���(OjDԄS��y�r^�������҆�5���A"�8�<zl�]��H�k	��n"�?�*#1c�`4@g�����x��K����+%Ⅴ�m��m��k�'�I]�v@�Q�Ȝy᎗���j�h��z��Ǿя'2 j�^��B��8}�u��������z �����r��z�0&�;Z:���v��ͳ��9�S���a�����!���3&1 _쑬�uuK����{��{ �Wz�i��+�"nҌK3���(h�>-�ѓM�����>��Ϝ�Ŵ�5�S(� y��\Zˀ��4�ݔ��7��-�"&�0�:_a���
���%�3������߄�b�2����b[��f0-�w�UMBcj��u�T�83>�8�Kq		�Р-Y��)�����B��E��Ϥ�+>�7GnM�����f�F�2��E+c��I����?���o�=���_�*>۔j�K\�����rX/��nSDq����r
0�������X�|����)�G�rg�k��C�M�Z`�����+�(�4Ba@ 
a��D����^�SQ�C8Ib�o6�؇��EH�Վ�?��s<��J_G��07�����Q��������x��͸��mA���>�Z��?-7�����)�)�����H���RmY[d���
�O��iE�'� -;�����[��7#|�{��5_S��z^U���>�6�A�μ`��?W�94�6D�g7������2Yѩ�F���&"�oB�?�eDTV�kW:8�\�:<��pވ���]Թ��um��bk��:/\Z���^��-���@ `��_67���=^g�5���Ω!t�M�,$��/�y�)�$��ʪ�΁CLS2��YXxo���1���^zhQ>B��%of&
d5�@"k�9����ı �1*x�_v�i�^��G����`�*e-����(T�mu�%I�q92%���L��ok�j��6�!�n'1&�}O�#��N��+lT���D�n��_�3�(��t��%�}8_�/�2�ɑbD��Շѷ�=zM2�}cU�?��:f��t9� �qׯT
����
�U@����[��< ]�g�-�ܻt-_���/��fE�f`Si4#HI'�p,^7� �{L�-ˢp��䱏s]
��K>�L�A�d�ݿ�x��~E/e�t��d�~��E@a��0`e}^H�&Y�G7����V ��1�Aʲ�k���<}��jȶE��t�0el��6�X�<Y'?��lt(\�K.��f��n���	/!�/#]��1	�r�����l��M'O0���#a��t��4#��ki����]=r�U�S�&�%2����6i��+ܮŖ�.M��!�;`���&t�������$�΢F\W��;h�>hFNvsB/6�D$�~ػ��Q�W�<:
��X�]�k($qr�����q"�L� �l<ٗE����mяu�	Z�w.�⨯����6Ykm3N3�/^⺇�n0��us6�u�A"��*���[t\`C�S�ӽ7FУ8�E�G�����SA��rͬ �-��Q���)5�Dj:���~�'�7 �n�K����~ wu�-�; �GQjR�����pYќe� 4ZXZY���������r:s)�z���C ���v�G�P�U�����^ԟ�op=���H�҇�{�ϪG�a?���A��G,��9W=(�`�����,Y)r��qo��^	0,�=�4f����?b�ַ�v��� �^��"���gW���;U�m�CI�8^  ��|_.�D,�~�$niV�������dv�Q��ȉ>lW7t"����`!��`.xo�z~]���܈���̞ �7�4�\*����� �0�2����>Ă�j�?�a��S��*�5sѣ�2�}�kG���~�i�����]k]"�uY*�������E)ҷ��+�nT�Ќ�ɒ�`Fb��d�k�KR��-S�n\�3,�b�E`��d@��c}>'�)w��t�-�@��b~Xv��j��c0��ށw-W7��+��G�L�����o��Hڷ��sF��1�L����p���Wql����}K�F?�tLS�@R��X�4qϜ�\6{��N�	n`�~ 1�/�7�!��ԅu��V�!�59Z)=*~������#���+}J^' ��?"?���rgO���z��B������T��^k���!��1I�ݳ���~7a.?�\g�Y���s��d�����Gm�=ZL��Fa� ���E	��"tl6 ���ܰ����Hx�	R�ū�N��D��C����W��l�� V0l��ۂ��#���k�L��ܛ�>m$���ڗ��hr��q���W����:6�DTI!�L�6͎�x=t���&��dĦT>,�&d*u���!r[B�Ÿ7FN�!�"��A ��JtIx2G!A<���'�轲e)w��/W�c���=e_\��VU�퍧d!+
2�Ǿ�"�[bDw���Y+2v3JZ60^�:��G�~g�I�/����h�c*Ye�͞2����a���zh��|�����Hv����23V\M0�o�A�thLn�{�O��XsŇ�i�7���U�@0�.6��5lp3 ���Up�-�����w_�م͛eP� 	�a��ĖR�x��fn���g�+�
����b	�t���r�a�|h�} �`A��bj�῿��L��}��9��2���31��s��Aɕ�Ib8��$4��J��Fk�}4������(��0���i�)��,`��+n�:�*�~Ff�w��.a3�K'Z9���'��If�j�}�'"Z�b�xSM�����18����q��.���-?�P�vq5��Y����LK�+a-y/��F~���ǥj���d*�5v6������e9\^V�j��v�#|i*&l��\R��,��C S�id��:f����"��+�y��L��/���2��"�a�ց��v��i��A�zXw�_�i9@|��T���`C�Y����Ɏ{v�/g��#N�Y���f�	�A.���b�~��aLww"�;�wqg��=��;�b����]����[�2��o�?w��m.�2��^h�S�pA��q��_TF��.FJ`G���0�@7?����gj	-���8\Yܲ"�j��AB��Ҿj����%�Di�����}���^���c����=��[	~ҏH���>]^��k+�L�|$�V�xKƛ��k���|>��sh�я�s��� ��*���܎��k�|�h��xx.E.,Z
�������ي��e��5#Bi�e�u�9%mU�׉FG�,��>xTY��|,���,Q%����R��4���F�8Z�}��z}�9[�f��U�����Qa�	��\���������W�hͦ�dՔ߷s��}쿪%�NHK���C�\ �66�n"A��L����A�,J�vvXT���)t�>ATע�[��7�����.��H1��3I��-�MN��%���ʀ5��v/G���3��$�u��|I�֭�MJ3�t�S���v�p��Pru���HNl܋%����fʣ�g��)�+Ѣ����=U��U;��?!� �����لV)���>g������<Ԭ8$vzg f��+H�:��������� 
g��E̖}N�l~���g�"��σ������h�R.�XlxVHYEB    5914     f20$h�%�"�Dd�TF�׿C��U0���é[�w�3��=�;+O��&��DX��E������I2���5+�-�����H,߭���`�̗�)�E����Pt2D-C��s�f��Մ���
PpD�]�ғ7�ǣ���I�@ɬ��ls�-�m��`P5�"�V{N����nT)��ބ���^�MA��-���Y��hp/3�q<���mO�RB���JN�F3�<�u��K�z��>T,;�8�{���I�������C�4�W��@5�l�e��":�2�=x|��hJm��wZF��NCz(�,���Fڤs����C�z�w��9qzvu���i�_w���=S���9c|�������	6�S�48�Ooވ� �t,��lO�9��DM�r��9ɤ��Č$�i�����%��c��edn�)�K8�g��g�����[5�%�u�Ҍ�xH�=��:e��8ϩ�z�{�#��-I�MemQ�"��냔%����1o\�RcZ����hbѶ��P�¢���d����%IH�s��A����pf��8$����q%�ND�<[��+�������+���o�:�Uo���GI"�"E�R&�0�6{�����ߎ��cjE�Ƌ�L��z=����}Oi���1�g��7T ���7��)H�(�q	� �+5���џ���a�t�3�Z�uN�r���(n�/��<Z���ڼΧco���+:�[�@� b�m��a:�i{�8�$����*h��KP��i)Q3}�dNl�D;������X���ۻ��ꋛ�Q�n2��nq\�Џ�ާK�v
3��д�N�\���AslG�l6�Re�}F2"z(��ܞ�/�纄�������+�P�"����"3�:E�B�|1Y}�3nQ���u�g/b�x��|�$�36�Oڹ#��b�.�Y���
b^����N,Q%H���2��<��{��g��8��V���&"A��S��(�7��_S���v&��rK60���"�K�
�>���,	��~,�ނm74����'6���U)JȗT�J�x�Q�0I�c�B�������|'�:v�]��B��0����������nhJzP���#ɍ�C������شC��E)hjo�N��]�,>�����	�&�B$9ćAK`v�t�z���e|�5�����%x�-�i}"�9yMv��urf<jF�*�©Yh���9y�ib��܏c�/6 ��9M���Q!���1����d�'�'��x����9�Q�y�Z�AJ>��A9A�� N5 ���'BP�FێSG�*Ժ�4��ڀ��޽�6�^7=�y�e�
�;���z� ��"�����7�h��l�)���]���p�3�ЏP��,g����{}-�vyhT2�"��jl�O0� �k6/�5Ȥ����OX�A ���e�2/c���<&"�[BBI��hlFJxJ1�[yg����	�e,�!U�Y�6s�y{��Y9핦��e�KzC�kV�6��2G	���؇0����e�@r?�6!xE-�����=u>ﲞ}�����W��VH+2%R,b{���7� A����d���]��j���X�ի�Y�����c>.x����i��B���?���/���Clevfɼ��,�*��u��4o�d;H+B��a(��W�p�9͎�p��wP���)�i*5b�n�b��@�]�@��[d���E_e�kL�]�?��Y.~�D%-��;��`�x����h0l/�^Svj��L�ud9�3�1�w�j�uS�ȓ��,���1����]�[K��#+�D��k��h�?}��N��=.�ӹ�-�F#=c�Z��{���6� ��k�Ňـ�h���R7�ii ��ig�?%+���e�D{�����;����7�����|)C�B�.�v������%9>lD�G��(��*����t���%�7�t�*I=|���1��zx"��]�"6(>\T�LFkVœ�d�on9���A�%�{��ɐ���#V���V�f��1�1ؓ��NQCJ���xp��̟lX�@�~��zD�g���j�VK鸮��I��t8I�}ւX�p���V�(��s�l D�R&�ԉK�*ፏ�Zg��ד���d�e��AҾ����=̩d�c���}����X���0mei�0&u9pnX�y��?�&a�^��nj՛ȣ�}u]�5��Y���L�����B��r+JW<p�&X�0[�EGkk؄?��=FH�_��D0���$b�("' ��j�v��x`,����Tz�~��A)�]���k�y/�-�ۭ��1���A>��di`��es�-��^!�x��X��dЁ��&݄Ѯ�og�����Ă��}	�J�!��D�e�G~"[J0�~~�p��o��=8��;+<>�%UW�b`&�T��W:2�g"���9gi�g����r!j�%'�;[�	u�`Ôu�08@Y�� dʹ�}���WgӔ�����$���D\6I�2!��s��F�}���>t7�\�w��YQ(����u���|q*H�H���C!�F~���`-ܬ+W�(�k�4�w��!�5�b���'���
��mP��`$G���R}A�����@ޔ�Ê�?��>�4�<���A��6j7ؒ� G�C
I��>��繌�r��G�|���j�z	���*;H�#o��rnl�.}
<q�43k�yWr��A[�}4-��Ei����t/K�T�6���DXEܚ�o���H�J!�e�r>]�� ���N3�����T�:�d%Y�@�	\8��K�P��/*{YJ��!�  �V��K�C*�HѾ����GT�׍�����r������2����XW�e�>g{���ǟ����E��&��M��T�ת�OYz����kլ�}���3��P1$z����|�����=�߀ XMmwk�"�Ș�PW�S�܈>NZ��H���4���� Jr�_��p�/�fT������Mǡ�C��w_�E����L���p�r?���:���|����@�e�Y7� �y�7�8*S����a�4�%��mɇ;�.F9�+`9*��_�*�+��O�ϯ��b��˨Z\��6���	�
�m(�b�t�8�Q+��۾��������\l1=���b��`%��ȡj>���9a�:)Հ ��,�jN�^y��z����S��#Ƣƥ��|�����wN�+��\2�!�N�(NS�SY�$�

'-����-s�kkZ�$o��+����g���c_yq�������E�!eҘBH���g������Q��MR�~@V�憤�8e����Ⱥ5�Ά�jX/�B"Aǔ7�+�u�`�X i���̝�o1��3{�H�\��g�և�@ҷ.
&���X�iJ�ƴk�:}�v
+��:p���2���ɝ
��c�[�Gv�\�-�P�I�?�9����/��Jc�DX����$fʲ��R Nø�M�bǝlL�	~ԽU�<jq��&�|3W� 1���������H�ق
�Z8��h;�|s��ת��GN��ѵ3_
6&�Ka�d2�c�V.YI!W�m���.f�=gt�H�aa9Il��T���[�J�x��_���U�/P�X�\Hz��o.��]o��@�G�^��4�d�RP���1�����2 �Ǝ��k󣉀p�^t��H���ϖu0���婎R���G,<>ty�§����a`'�V
Cb��'������J(%2C�R�����;Ҩݔ\^�?��tpt���S+F�C�|�u�V�J�k�&���� �l