XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|*��t�P�H��y����A")P�0AT`#��=�ilS�w2��R	�*Znֿ���o4F�P���N�ni���0P{�D��eqG��=*4'@��p(��~���v�b�і# �Q��T��:%�
�lc^�i���vf�}����C%+Q{��l�� �*+z6ʾ�A�����j�1ŐB�(q۷̥.�{r:��z��~zX�E�"ٝ��vu��3 x�i�"��܎?��ㆧ8��Cا�_|�6E`CO|�D����(� %�lo���u^m��/b�ʨ����=O���HD��
Q`�^�N��Q�0�B��Ӓ����;]���i�\L����o#� V�� �`�HV����ʚa}n��S�3�ڈd{%���6��r�VW෥0[���g�����C�J�H`��HS3��%;�5O�l�n��a�2�q��:I������e��L���Tj|���k�c��P�Ə�o�AgH�X�=�����X��U��p�9��c���$mT�5���$�|�>��W���.y�'��m|i��/~xM/ԭ�Q��3Pb1&���,�����:J/_b?� 챁QL�:na�w�$�Y1�i(�J����>�_��.Ǵ�c3�L�UƢ 6�`覆�����yZ�fUʅ�0�ac+�0z64��iJ�����T��z�=�0�cx�`Q_�~�v�'X�"st��S����8m�5�E�,�9��M]:!B�v�.UXlxVHYEB    fa00    2260_�)>]_����������~t�;�Fp�|/ٜ��ih��ʹ�4I`�����|��b3r&���p���{�g�o�P 3g��js9�M��s&_�X*w���:����Ne�}�G��&��0S���	%�����渶"�E֑C5]#���U���	�0�6_�Z�j��(��#y��p�����:x=3h|ƅ��Gq5�:Ā,������4es<�����Yh��m�x��퐨� �_����v�.��r���M\�j�s��r��[�D*����c�����8�ը֑l�̜��i�!�%����<_�I/9(9.�����Wp�7Y6,�,U�z�~��)��	yi���4@q�9�f2=�՚�����~ya��f�$�Cq+�[O�9��C)�;�}Eֆ�wV���!L���E=��IU�^U���E��/ؑ�贈c������{����Uf�}��v�^��F¨������HIp9�oR���ou��J(> �ϟ���.�p��Qw�s�fY�l*W�-�b�O��q����A�����P�$�YB�9�@V୻�����.ڼ��g��=}]�}�s�G���(��e���������A��ժ�z�T���7������u(��a�c�s��b���$�8{u�����]<;A�3�XS�@�ewo7v��A�e�)V����Kʌ
��x�e�����0�Eq���wnB���۠����L�Z�QN,���)�c��Q�8rD�m�I
}D�N�ߊ>��0tbgSoc�D��/\��d�Bjvq]ܩ���sǭg�N��ɭ�r�G�L����oԴ��D�\,0��ܭ{7�����T@717�Pga�nx�{�_�7�}�B:�{�8�`�!YF����[$	$�g�?o^x�ŘrM�v-�y�FT�¶j�����#�ۙ��n��nA��e�iqX�K�w�Ɍ��������l���4�V]��3m�� �iC}�^�aTP��o�=X�� �[=T�wǘ1�y2��LlV����HmZ�X��%�kblXA�U+��u����c�n��mtH#�v�/S�Fy��|����cҗ@WEQ�2k5^� ��6���'�5Y;�+�"Dp/���7���0(vE��Usj����2�H�b)�VV��Ď��O�q����ΡH��a���c�G^.���^rf{�jZ-��D$��#����%+]�;ݩÔ���6����'���qJJ�-�Z�����z,Q�(��m�@ �+����=�Ȼ $�9�������ֱ��sд�w���?9>m�W\�b�}ͥ����6�0e��u�
���N��d�R���0�����nDv"E��`Fh�R�V[^�(�q5+���o��an���=B�K!�h�;-�D9G'H���˗㢶9����������j>
�pY��n9��U_Kّ~�!�Q�:�nZ�!x�O����#�V��.w�q���Z��_q:�:��U�|��K�gBk=i!�KO 9-�4hj�r~r/����p[y�( ] F��v��rA�ġf�z���
���Ͼ��ɂ6�*d��C<_����e~'�T��bo����01�2�+�+�R����:���� z��;�'���}�\�^�i'둂q�2���L���q��@6%��eoz��Ɨ�~(��Gu��/�&IZ��SU�1���T7%�,F픡�٪���1������1�aT~��z�ln0����}wƬe�9bsx�}��š`��kۑ�'��P����52Ǐ�y|>8�dH�h�GUz+d՞:�a&n�vYl�N����z��;���:�p(.�;	{���7E|�0��AF��O4$VX�I�u	&C�K!�:=yMf�G���7p��X㩁j&D����d��9�8y�u6@la��<wi�Ϯy��Kv�*��\�&�L~y[��(�i���?6:��AZ
�	�A z��.:��;�n����@��ԏqV;�mnK5@�\��#}�4�rmz`��Jl�c�g�$�m��[5`xa�Ě���T���#r_��o&�=�'N��������K���L��)1�=���C��m�_@�ፇ�@�IڦLWEl�[K�É�Cϖ�i�#/�c��e�*7m�Eڱz8ü���{7ߖ��!��jG�p6y�pÿ[��y�<�a�Uέ1-�3m�y�M��s�8�F�D���E��H���P������0�
/�P�m-o5~ϫoh�x5A��0�W?�:�a�^bV����>�Z�{� �r� ��迵�����i�}s!���M�򏤱�������)eC��RY}��LQC%�I�h�K�˽�;�Q[�Ui7�{�w�sJ+r���\a���{G�6��S��q�؜��cc���6�A(ZDVyL(q��I�}�(�T��Le`k�ʇE�����y,�:X��;�FT�p����z����gR��5kP���U�ڇ[���������1%F��/���d\��ړ^���u\.�>����S�7ٹ���Y��������]Kgh���Z�d=v|�{_�v��	=+o�e�cC�Fz�$�D�1��%J%|�������۞�}mo�WH=����p7ƅ}9m��
hK�0>4� ��m�(^�u��Ԝ���zzT?��l�|S���At��@�lv?�E^f/)>c����kG�����+Y�e��=�¿�~������C�}h�	7��5t_R��(!�1����(|�R����hKWyZ�=�e�J���!�i��p�d�k%>�n��E��ҍ_�j�Y+��i�'�jy��B�=})XU2?ɲ"L�;�k�D��>R�
��P��w|�����4�^w�+9�jɜ���^8��z������E�� ���#Bi�$&�UI��#�c��|��:�M�S��o���u�&;f� � ���V����'S��{c��Y�=?yr��Fx^�r�T��8�`ݥZ�U7&��g(��U!���-�*�����{M��ʿm������w6�@� �K˵�"��#`?��P��[�4jR�zl���9����pn-]�́���4͓����jD����:\���	�$}9�����m�?,���5�:rE�2@������ [>z�CW�U]�3&�,����H�,PZ`�z���Vl~�0�2*y�]�m<����-��e�]�Y�ۉ<y�?���Շ��Xk�3���PTj��#�=9�������r��+�y��*�t4��ö,�ꤐ�GӍ���	�������:��ۨl+0�����ȀcH���5]a���{��_�;'~�����p9vW�A��z)Q-���_+T�����^K�H��p�`N縪Z����R&�e�uϔi�1��gʍaO��>�}_���������yyH���Nړ�`C|*����-�p3�C�{�;�5z�Vh�n����є3�����3�>!5l�5�{f?$�*$
k�����Q+�kG���;u-�y�����n�Ƶωښ��Y��P�O�ZJ橾��&�L����~��.S<�T_���W��B���C�,�7|Ȕ:�Qm-)���:��a��.��1�|͢�2Y�ѻ�2/���������VB�E��q��^���rɪ�b����P��r�{}�,`����,p���x?���1=m98��@mh�����T�8�9J�ZC~ў� ,�ݘ*�+��/��3Q�h2�Ds��)0� ��7��	��sE�(��9���`�W�u.���Bsda��ަ/!.MA�1�,�����8^R�|va�"Q2�ǿڲ��LJچ�ZjȘ��$.�Ͱ��|���ǧ�]��X$А����O�;>���n���"�����ՏG�����z\�
�w��]	_<w�El��-��@��'�szd|+��}�8�P��g>�jc@�P�ư��,9�7/�7��d�*S��P����_�}�Bp(�ƥQ8�$��yB2Z���a��Z�-����+�iV�uGp�_Fj%ԼWkK���ȈE�jT���p���Zqơ�,��(>�n��6\������B������;��Ty�hS����/n�W�:0���~}~+�̡MAѶ�Nw���L��:%�b�����C��JG��z����|	'��!�N�������4)a���0�k�J�_��0��B����
�0�%��ę���q����,S��X���*	/9@���kӵ O������b��`��b�c���S�vy��b�G�{�{|`^6����Z
&̵j���P��-�5�y����(�\�A����;�16֗�sp�@�g>eN�$�>p�> �m3	}��m?S^�C����	�`f&B��H�I��s9vS�(�"��2t���7��d����ExZ7�t~o�jR��7+!�1�Bǋ�'���+ˊ.��R���P��ŸgXn.�JI�ԧ wͻc��y��Z
P^|��q?�,�𴙀���~"4�݄��}�J1���#��573����("�@��wj9a���ᬏ�m_��WN�Kt�gM�:X��D�� a4q��C�o�פߛ���@���KA0^�gG���VSȏ�(���t�ʬ��duV�������+w�\-�|������b��dWO����8���+��;V{�.�.爷�U�"�㚏�F�u�/T���0�$	8�E�v;��a�h��\	Q�]��)����s�^7bO �?*l���#���FP�ΪH�ev�;��_�&�b|2l9#P�Ift�"'=pG�fȻnˣ"
�6Ͽ�wc7D� ���
p&��m���n	�d|�G_��>Bч�2�cg�R���I�?��G�O?�Խ��M��e��ֲ/t��:��ߴ�2QE�u�'3Y�ֈ�&���u1v�o-�.��.�{�TK��H�����XB�8y�'�JFX�ܸ�UA�9�Ԓ[3�[�������oD�����2S[v�V.�����¥&�P$\`L{,������>,BT�}��7|;�+Cj0g�J{=6�h`�G�p֫�
�;�A�tߺ�ޒQ[F�@��>]0�l��m�p�]D:�������t�$����j7J�Î�����ݍ�Gzs�!��ԕ%���~��i=�p�$ވ��`M��٧v�.�m���aZ �lz3ڷKe��(�K��)���9a$)�1����u0
�Ej�-/�H�+������"*#��84
H�d�
�����'+�hMz?���n,�5M5�|��n��ëw��ɨ��	%A���b�J{�zr7(��� ���N����=�utu�վݬ3�̆�SF��x�l�k9%u�i.@?N[aw���r�{�|~����6�pp@�;�&�Q:�"<�7���cY%#e�w��us�Ԃ��l�hq%���&��|a��lNNI�Y�u}��|��	M���eL�ع�`@�=�OAD"
�&���2�+Ӓp�5~d��B�*H�(_dѡS���3��S�8��w�X�?����z�߂Y��[
R+XK�i*Xm���~�`��u�N�ez����M8$������>���4��^fo�<(5I��V7�}uE��9jc(f�����k��4n?s?��1�Cm��*������Oˆ��J�'�	P �H�� �eB��y 6�*?�����h���8y'�4Դ�R"��L�;Y�{��=�V_�	�ԅ�*cb�1����L���p1pe�}�m����:y��²T10���ډ��u�p���m�<e����I�-_�9̸����~j���8_,ڬ��Zy���������@*?"Q�]Y���9�*�d����p*u���<󬚰��J�y��|8�G��57Bj��?�ҙ:�"x�q�mN����#�逷���qQ�`��j�$��+�n��Z�0�3�_����Bc��C��0D���^jtcd�E0RA�<T> ߣM,�iD�1�Eb��U��x����O'� ��X���G2���쭜��@)-�����Z@-�B��=z��f�µ�a��.e���Eo?�Gc�vP�6�M�)�d�P����{*oP��{x/�'��@މ��j_?�-4ml�?f������<G����e�⠳;}�4`�M/4b�H�r�"��^�f �d��p�$\�����ufY�@��Mַ�K�7�M�ᷚ ��SY�"�Ň8'�)���7��1�s�od�p�'z��L�	��M8����2]��P^���ն���d�9��U����h��J�P�Qؔ���sF�0�[W�o���jk��H4=��8����>�*�z��ej$Hh�#�ľ�%�P���HT�Q��g��3?���$�-�K�	~R��U'��yP6�Ş�/�Ȍ�O��Ec�hlɨ\|ܤ-Ѫ0x�Jxap��͙�.cf�mhk�5*C����˳
�M�*`����B�\Ȧ�Iw��d��	ea4�#J�cG�N�7KnsF0#�[���L�I��g%L;��hH��o `{'"s�8M�A�:!�:)�Qh�����)�{��d;�9: i[7(��x�Vx��+�4̎ix^�F���)�� �o01i+u�"�]0�����dU�`^.�O<v,�������������S��m��\/�=[9E�`��+�7GRh֘�
]PfqzB �Y�_��	K.��Q)GB�$�/%�rmж�Ί7�v��h�6R	��ZGM�v�ɏ
��c�}A<�r�+d[}��?V�)�I��U�:هvf<�Ҷ�G
���U�U�R�_�ۿ�7� ��n=3Of#�|tIj^��h����͖j��u"Q�
9v�v��l$7�KDy�4qN��Ƅ�+��<�5�}�>����;p�z��L5�ݙW4d91����$ +�ߚu�ξqlm���c�'��G�/j14�Ju��`�'z�eHl�"��V^f�$��v_�9�c����N���P
����L-�3��`����Xul ��q����R4���P�)�8A�5�"^S2z��� .{��ڛ�][��Fƹ�Յ�l-uFh=jF���v��"G�)��e;�M/��{̤��B ������r�]���dəF�S��3o������+�!���������CM^���&Gܕ��w1/F9ܸn	���WHCt3�`Y�������GS�M\r����*e�v4�D��2�+]O�\'��X�^ �C��4F��0i�'�R��X{�Q�]}��z����TPk�)��pțH�{��z���%�ʥ_��+z��"����eR��4���.u�Olg��\���s`*�nZ�K��5WƑ�A�{� ��;� �'��q�q�i����6�/�+_Kf)f��當��[Jf��?K�~h#��B�ߺ���
�v�%����O�b!g�H�Z�*�Ӧ���WE�/y��*yRDb��@L֞9yr�Mu���Oe��C�ʮ;F�p9 .���uk��~�n�(6�s-}z����$�2 ��"*��	>��Abj��W�
'H�չ\�ҹ?tp�Κ�yQ�����׏
����/hhn'�p�j�&�l����@���-�� �Pr��y)�eh�K��<D��ms?ƭ)�ز�r���:��HM�a�V��ԅ-�ކx�ى//A��P@�B��r�t�!0��.(+��)UA �~U��9,�4r���HG�W�+���=V���Ԉ�v�/�_\a���3�Z �%�w�{�S�`� � �����dc���	3ע�����F7�qUG�WT<��}��֔<\n9���Dz�g��ь���X�v���Xb������d�
�*�0��k�"l�s29���O߼ɼ�z���y)e^�z-$Y���&�m�e�곥��+��ޣ@m>�=S:n�EiK���M�9���8٫�~Ѽ���~�����X �"�(+���=�"$?�r��`�M��7u�5M�Q�n��i�C� 5�����]�׏`�iJS°�@PK���� roO�:����G�u�F̢jK�P4ȕ�Iu��#���x%7�U�8iq�~�4}EB	�m���HZh�:�K���|���T?�|��׼*dhk[s��]��
{T_ZG�~�B5��R ԋ�}]�jM԰��[>�˵�23�����_�B(���!���6�t��4��(�$�V%�q*@�<�ͪ_��K�ц����]|��/���d���L87�!�PӉN@���"Hy�\����ݲ��O����g���狫�~H���  ���J�Ƞ*n�w��s�!�V��Q0��em)m��+�͊���%��I��z+]iYxt��n�@����;��*\q8Q�I7�\�7:ݟ�t<1X�� �t��nhI{)�:����W�Y���T��=���e	5�FB�V�{��~@q�(L�z��Y���N�����#n��~�ݔ]��`Ŵ�8]a���ui0�8�9�6P�{���W��v��~��&n/J�����y�K��K:����%�2�FM�s͠\�h��� &p�-&�*����jV=�טsRv���VC��;4�,g��i����O��t��n���SN'�^I'��5��t��"�$k� �Ɔ |�j�9[����%Ɯh��rk���F�$��!V�=��	�8SU�ݭ̂i>�ϓ{������lr���7%;��e�������N��[�Yv��1H�x��<��jWX��o�!�XlxVHYEB    674c     5c0�"�ƷsL��3Y'��F�1m4G֙O�����)V���0���l��_�����ի��
���d|��:N�h^ŲWo%�#�ZC;¿/ߢoh���S��b���e����a+� )�k�98���,��G4r��	�"	�N��8Ϸ�'Q\3��1'2U1�k��B�`Ds���w��3�΋����9A�,�qF�h�n>8���9�[��_|hl/�����3�/6��?�{ �[��V#`�j���G3��yS&X$��-1? L��G�`&`�-�,8��QC	<\&�J��Z$�%�dڣXJ���w������%��j#c�^ �X�
�.7<��V��>����ʴ���c�t\��BPE`�N��N�N��N�uF-x&��n��V~*�ԫ��X?G�O�u�$Ѷn�`	������PY8a����R��u���{U�x��x��鿔Qq��ś����ύN�(�XOfg��=��>� k�Uε���"����ժK�C�(_	���L*/�U=MVŒ�u���Q{W�?��q3\c�g���6rȮ�(R}��1lF���K���'�m'qs�f?��[ɫERKOS'f�V[b�K�+���D����O`��bҜ��� +~�s[����;�bOG2�������
�j���j���v��o;�`g �^C����C����{Cv�_p��R�R�Vq�b�ؔ&֭ٙ��iz�b��-b�9��w1�5>Y��!_�}��YQ��e*=���b^䱱^9���9�Y��\?���u$��Ύ � m��l3�J��EE��y,���%�M� c�(��H�W��;0�J$t����˫�7�A��������:�i#����~����C^0 � ���ʃR�)��8N� �hRR���k��*ƪ���i4y?$� �9ɐq^�[ż C@+.}7FR�:ׇ ��Ӻk��5ȳ�Y右Me>I$�@�˾\Hs�~�ȣp�|ײ����nr�k����{���Ưp�W]��ɱ�&T�ltn��X����%S]J����|#L̔6�n��b1�)@��9ƨWl�A;Gl�#��h[�U� 0Pe�S���1C�Ǧo"�s�p��Q�*�_���[�.��۰1�so��� �.0��5�!U�Zv����=� ����O���By>܅��z�fĢ���p�lx4G��U�͉��q�����nƳ8�I7i�x��T�/+���VoU�r��G^��~�*����ʳ�!	f�Ɠ]����5�u
֧`"�ة�u.:J��&r���ˑ�b2l@r���l�S�r��4{�p��S�GWA��G�1��<�M {�Zw�p�
"�g���#�{���mȨr`�S�m���߼�-̮�h�r�)������en��U�j��#뼚ъ�s���X`�V���]�ʢ��t�U	�1�\$y�-Eye�Q