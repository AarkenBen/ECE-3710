XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Z;�/P���Q���-���観ZY��,>T���z�d�b�_Đ��/"�ܻz�%�k*����6��V�5V��	&���Zӏ9�n����/5�+��/��dnГ;����z�9�f��b��V���mT!��,,����a�`��%=��C6j��4#��?%:P��X���Y��T�F���T�[��{�@�Sy��;12EvI�J`<|3���0��@61�d�Z��Bl�������V	7��R�ƩPF~�l����Q)��h�-/��[p�Zէ�D 1�5��劎�Wx��	�>�������"�nTK�,A{%;�"D����l��mF�lkC�d�L�kU��M��ŉ��6*�./q$]�(qOĊn�P��⋛WC�lu%;�$�C�RBJ������
�r�w[�/y��y����0}7t�o$Z�)V��T��V�Ӛ�;�plݎ;�u��#�q��+��]���Ӕ��<=s�ze [���-8Mn'���3)�)/�M��C�"�&�#�^�`a{�f�d� zNO���y�^���#��	�1����S�t�U����5���%�{��2���t9����
}d��m[d�B�6V�>-�����Hkzg���e��8p��:��F�j~��4`���ܟV�����ar�qb�`�	�O�вs|�B�Ax�i�i�����MS��f�Y��z�d!�·U>kL�]JWK~P�I,��`�I@$AK���^��*>*�XlxVHYEB    b631    1a00���&q.��̤�p;�$D�R	g`ݔ0�����L��:��}�woإ�c��fMR9y~�_�x���I>3ˇ���zC�y_j��V}]���CJ?S�8��9f�,>���*v~Ѫ�r�!)�wnݍ�>��BN{�:��0�bu��P�54J��]�Jd)���נ`��FV�I>M��)�ƦNi�ˌ-��	�Dn��渜Ŕ}�g���^�V��詮f�-��]�0P<6	���a�� uŪ%��5�~��	�����I��/�Z�2,��U`��$�~Pxs�h[��Z�Ͼ��Ō�0x5Ks��n�΢�O���Y(����"xwD�P�h 4�&����<2F���\E?cCv��� �����Ț~��4u/Å�!Ƙ��:��l�y&W=b���b�C�F����t�ڴR9����Jp���Q�S�I%�$Y4�����������j/����m����E^2�l� ��1�t����S�'��ȃ����}(�3�%Ftw�������5�����ն-߇��fR�{�'[��2�a�*H��+I�H��=C-�9��0�ˏC��J�&��ưkG>N�	o�li?����V�Qrd���<c�hzT��x߅0n쌔3�`�0�!ɩ��Z�PƱ��k�
ƀ^�#g�6e][�4R9���A�*㕂�09�y���N&~R�(o�.�.E+~,�Ꚓ�>T�M�:ST* }(��>��Z��,c�?|��x
˲��g�~6p���}i��U�H��B�wd"�l7����6���kSތ*+�����X��[L�#��?�ʆ��ɻ.
+C���E�Q^x�{���Iu�~ N��}Z�LJ�s��Q�-0���xPAon�5��R�*\5e���Nl�HE~��ku\x�d��pv��"��o!]M&2����%)�1zR�#确��3�N�����2�c��V����і���>�ؤ��8��C&��4��{��6���pG��!����n�+/����z����ӟb������s�+@ԑ����ɮ�<��� �!��K�a��>q-���H"�lD�������8���(f��2�=�5;ƺ�b�̃
�l��Hcˢ��d�2%�/,@�P�@p�=9�k� �l���y~�g �5�Y���>�3`����yV���샴��8����T���9�c��P�%��E��t~����/�^T���$!�K��DO�a����`-ܶ�E����G�f�Z����RZ:��^ 6|A#��m��M�@3y�-.>��Rn�\U���J�!�Ci����o��l~��k��|W���c\}@�!%��yq��(TS�Q���2���.ᄊ.kZk�fߧ��)K���5�v���!6��au��>�8f���󛰡i�3#��&d�ie����3|�})C����< u�B	G@�a��gĹnr�)�����)��A�9ψu����ז�>Iz�r-��}���a�����́��3�`���PN>U.Vh��[ȍ�)16a����Š׭�������R����fr�>!V<���ײ.�^�sm�� O(Z+�����������4�����,�"�PTi��o0��΄��8O�ۮ��_۪�#}7�������`��Ba�ԋ����y	���J�8xk��C�W�)H?B���Y�!k�kFO�M.W�.��/�EXW��y����Dk���wDO���ׂމԡ���B�����G&F;�T_֥�{��ѡ���sJD�7��3�{7�q�,�pҐ��D>��+���i�w�Б�ȅ��LB|��E��R<�/O����2�3b]����;"{���f tvcs�U�0�pΖfY��p,s��s�ވeh-:z�L�j
 ��~Pg����pY��6$�B�����G��	6.�J����P�S��;��Fo�Z����_/ a�%]�X��6?]�Y�!w�;�;Nr4�XIֽE�&2��MW�}Q}�n=Ws%Y�S�7�� f5jg��X@|�� �Y�f��a3?L�u
��U�2s�qCǖ�8��yΙ-�eM�?���A��4|'XL_g{���t�tZ)S���E����WCP�� @xG{.3�UH����_��xj_���U��!���\�tc����F箈!��Ă�іV�<�u�N(�$Z&z�|a¹��hy�w�"R�B%�	YO�kU�`B��ǰ6���f=�0��8XoK�ճKhעI��z�5���;��U��v�Ry	ֿM�_�c��6�TX�t�᮵���ei����������!T̹�%09���|f�x�U;�L�8��L	(&/<��1��G]��N�tv��(�t�8�W������
�R�2�6�u0ĂuD��>Z�x6�*P�W(g*�&�����n�ʳ�:�
IRr�_���[�z�oC�mA����l�6�u~(	1(O�����AE���!� ̩/5��u�������B���+ 5����
ȳc.�21Z!=̖�@�����x�Or������BYPn��� %���L׌�ZwGQ2Z&g����E�:�'��0�	r����N.`nf�Yg͘G�T|�Y���!�p�ѧ�!�[�o�C��=��)�BQ:�	���[Gt�Ν<GZ�la�;	փ�ҴB���{Dt�w�H���D6^���m����:)��D���<Կ�B�s)D_�A��K��<Ű��dS�!�ƕ��=7��u����!�<h_��<	W�g�s-��ѥ�ۮv����oݵ��H�A��x�����G��2|�T��4k�:o���,��9�U���7�
��E2�
5��i����D��z��PRȰfz�lwj�-@'��'@�ٔ�E�������
7)��M�2�'}�I�d,��\�p�ݚ�F������wZ�d�P�i�N�Noz��mEl ��֦�� ���h��k�8�>X�L�{�FUٚ�s� W7o���&��z.�T��<!e��b���L��s�е7L������紉�����ܔ��B<�4�߿�܌5�q�"�awd'�mBgM�$EYB���MI�~ xьܦ1d�]3�dp�+�A�>*���7�!��n����V$��)�^}�)c}�����Uˡ��1@�xh#��t�S���} q;�,�⃂�ڹ�q.*|���k�%���:U�!���h^P�iW�3���,��l%w�0-�,>e3�j�����؍}�وȴУ^�C i] }�_�3B���Ԥ��ծ|[r����3���c�53F�#��3G�	2��cle �aǿ �nx]����G�,II�U1d�����Q/t�B�]u�H�� �3^{��b
6
+��vf�;l�V�YX`�|�ݡ璣��=�*3��$h�=��TxFN!܊��|�ѯK�/U[�k`�7�1��''�yD�'�˟��Bc:���A�=t V|v]��Eaj��ʞ��eT��LFTD���96��O�i2.�FG�Wd;9vuuˈ>/�\{���F��*)�W(&!\�ZHx�dQ~~���1�p������|�_T_T��İ�2Z΍���>4>�+j�I������ُ�������C�l��;_:A��u[� �A?`\�ҡ\)���:�=���!��+���F�[U�ȸ���;��s�<��31�6�y
����v���üRK�B�5�vg�J%����ՀC:b�U�&� �*�N~�[$fC�+_������mgz�}�[��eZ�+3�p՚j:�*n,[ay�g�k H}��u����v�ش�d)V�k�b���+�O���S,��� 7c��9V��ǝ�G �&l�wY�r������@�n�d��� �r��F�Y/�i[��f9)m&���f���? ��nz��F��3k[&>�9T�O�4�	��9��h"��8���iԘ<�(/�^�(�}.hc{$l�;8��Ȉ��g��Qy�xC�I�/����]q�h�Ϣ��z��э�����w|���L�"�H	��5�!�`-�|��OX�9vP\i�.�˂�7Tg"���ɰ�=6�� ���Dh_���櫶�삲RV*�V�I@���C��J}j�!�x��߸��n��sG�s��m���C $R�<�b��Y�c��}����#2
d2�07G@�D����H�GT^�` ����5�iw����V�v�SVF� P��KE�؄�=~Bk���U0o�$e[��G�늹b>���-�#�B%��r8��Hw���#��C�2Ⱦ����y���@���X������&O���#�^�4�y|�_��q�W:����$�Q���j��)�e�H��]�,�>d��|�p<4vk� ���2 ��H���Y6�����k+�y\i��f�������Tk�*�6{�y�W����O��8eO�@����F�{�]:�7=/�Zes}�B�϶��� w�� `ӡ�%����0֬�Zj��w�3Z��fncD�H�γ�u�I�����xMG��&�ݝ�Z����>�KE�Ph�uF/l0����`���(�T���gj� P�~v����r{MJ��f1B
�:�>�`����Hu}����fK/���NO�`���}�{3p	o�b�`'Ȣ���X�mRnv�#{;�A����6�~����Q�gt 	3�0����Iq���>�BG_);�c0�PΚ�CR ���4���{�ԑ-P��H�e�f�C��q`r��Pas��f�	ԟ�l����8�-_�-[6�2��,7��,���ł�,ԯ�У�I�>��(�f3�#�FL*���H&Dх�޺8�p�\�1=�}��X�����٠�f�����|�ˆ� oQL�(?|{������M8�8�*1Z�A�J���;:V(w������r�1d$4��a�e�ˡ8/�$��L8��PX��}�,h�B���u�L��a��܋=&@y�?�,ӿ���U�U|P{���
O:W����S�D�k�t8ʨNhfĭ1z��dO����n����bmP(R��y��Up6��HMx���@Y���M
��D�{�T0Ҙ
��O# ��Ԝ=�*.��{�M�>I�����F�wgLF�����
HG2Z�KrP?l��d�T<(T ��یA�6s?%|�� >n�g�8LE���DXGXEm�ڂ����ȉ�£�v��V��x���m�s�;*�����J��-)3�{҆gh�j	ޫj�.������78����Ţ�<�N�� e��T��G<w�rS��}��f:��n�sc�΃����ӕ��jB��T2���`=�*���	����܈�w)�؟Ot(^�3����|k��SA&�H`����ħx�e)M�RN��Y��A�^frV�a<� ��V!��7mT9�ao�j����y�������B�^�[�8���_��]�&�v��`(֒
:"g,�+a�
��&� ���`i�rL���x$xc�'u�po�v�=�+�) l�߃C3@�^�,*/Չ�<���N���`��F\�����6�erk�A|����F��a*��)ys������B�/�]�M�b�r{Զ�WU<~�Yh<�Z	4�ꮇ���V�|��@�R24Oz�L���ή�i�R����1!�=�Yb��wƣ�.Ӗ����� 6v��h���4��q?j���.m�j�ɸ�D���`���������:7����7�>�P���Wk`��_׋f�q�>7 ��7{��X�FY�X�I�~�Ë��T���ۋ�țk� ��b��x�V n��Q#ţ<��Cۑi^�$�.�.�	�K�(<N/$Ȟ�/�Fcu/��F@#�/Ł�B~NW��"��u�w�#�(��ӵL�2|>2s�mR�ky�Dk�ǈ���.3�Nď�Wƃ�`�=�w�$in"F��J#�g�7VM.�}H�l���dt���Ϸ"@���(����\jy����7:!���E$�Қ��Cɏ�+�/�y&~������H�o�i�;�g�p�Y��T�7�ʖ�=�YTW��,GB�+���3E�h���F@�uKbP�iYth���c�Y9�L�J���.�|�]e���z�x�Cq*��ڮ��s|[~I�S�Ųwp~H��� ����k)��}{�)7}x�j`����Ks��"�=�����8��Z���ub�宏��N�QL8]Q�bmaT}6���X!P�ifS�Yݭ�l���O0���nJ��q�S��%�l���8��ϱ�H��H���z�D�6uD#xuCSu��>Z�{��ƗjY�@H�&��i-	���)qv��P �F��0<�E-��=�L��G�����5~li	�Y�%����}��/�}���#���ay\�9��� ����,'Rc�R��]:U|d�ߟ����\{ޤ�����6)�w�Zz���veJ��/�u�e:26JE���K�O���U����\��Ͳ"n	Ib�4�g� �l�[v*�����4���*����V�o`A]'�P{�FvJ�kE�ԑ�Uo��Tso���]�6�,NVRA��K�LC]w������s��^.]J�����̴�