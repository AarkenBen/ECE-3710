XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4b4�L��	�E����_�*+RLM�{{����4��Ĳ�v1/g�~V`CcX�j���������r���֥�'L~e:n"35��	u��/���+�W�KQC��~7��X�I�Q�{(�i�9��x�!DUEՔ�p�`ۂ�t(�O�o� `ц��*6����lF���fN[��� vO��y��+e�?�B�v��?�^*�D �6}�_���S���8�w�(N����#H���1ϛ[�4VdG�˽;��gx[�����ý�'1���R�v-�4���6�\Nm�DJ�"�)�]Z������b+�l/��|��oB��T2s�-����ϰhm�n��.�?�+=�r��,�~�t���q#�1�IAڳ���&��ԋP,���'Ab�d����X^B������(�g\�n����E+��R������ D�R�/�k]lR������N���B;���P5�ؓ�q䫺-ZҸ󾫌#=U/h(��y�n���-�5;`껷��DrX�8ę�c~��[L��ϙ��-�{E��Z�r[�J��(����><x/�r�Q�z���R���<�ez��i;��l���I��=�$qNK^Rr>�O�����)	LV��[�o/Й���Kd�/p�/�W���;j��z���<7z�Z��ir�"1bW!H��.������;�n] t6�zg)�)M��Mb��%o1>>Z�6h`8��n���Q��O�˾ �#&�fP��7���h�m{o�XlxVHYEB    ea93    1880l�[����=U�~�[J$%����6Uwm�\�f�5�!2��ř�xxΣBD��Yz�w:A�-(B3���K���N����l�~Q�u���^jk0��vy/C#U)p�I��ui:K�}�NF_#I�jʕY��eD�, R#�b-W�&�ƪN
�̗��p�˹����6����Y����uO�K�x؉/�"�`K�"���%e���E�E��ިK������+��'�k��t�F�o�d��Ziw�����nt+������:;o�N� x��[,��̐����,�W�FD#ɵ1q}֧xW��z8,�����ԫ�c<w��x�Y߲U�-�嘇sbWK74�RM�6ӳ!�}m)ͦ�s���m�%Lu"/����S��T�tƂ�d/�5��pN�!G~$XR��t�sU���<MZ�p���
���o.$&h����.��6g�`��sv���N���ި���Z,6a鿎��M�_Y����Af�*�N�B��n�}��;ޑ��굋���ڽ*��И�k�����
�9z���SP+��Ⱥk�	`;?�i԰�Vw�&d�r��``{�Ȃ�b~�Y�<u�59�\�H�����GF�Jx]�#l*��K+M|:���?'�������e�'W��M1��í�~A��EFeܾ�b��?�I��w��@0#χ#��6&f�N2���k,�0g/4�.��aQ{��C�6��ވ�̃��PĂ*9�k�Ԓ��@�XW�����Tf�
l�X�e�"��)���x��p���$��$����� �[��PjfD�l&3oQ7�I�\�sh���~��H���̪*���11G�7�f��<��X@iW(/��Bq�f���Է�9���1s%t�/5g5�$qh�q�?�˒�F`~��G���	��bq���x.kIhQ_5]�,�X>���w��8�Mn�����q"�&v7}|b-�K���~�����1r���1D;L���)����x].�^9	&���9��k�J��.����5ޚ'c2�q�l�77��m�Q���bj�`��y�	��}XP��˼@y�����'u�7�K�ז��ֳ^�l9%����Y/�����OȕuW\T�	���~�l�5����i�^�]�Z�)��IAֱ5�#~r�H���&�Z��VP}��{X��},M5�����ߑ
��|����</�_�ք3�lU�˥+6��"�wa$l�J#XV��挋/,�M=��*�ă�K}����f��EXGhA�Fh�u���Ycϣ
>�O���j�ԝ�,�N���6�R"���/�7r�'���Fʰ0`�ʷ�o�j��X"T�n����·0C�ͥ ���:��=����wQ�����;�z
�����P�i>#tT%�!4-��.w�X�D(p Y�q%��v��:q6Z�k�\�ۨ�(%�c����yA��+1[�MT�7�ͬ4�'���^^�K�4�i���8�,T-,�n���y���5X�,	��ʐA� 
^�o���w�L}DC}��T�X������@�rC������LAd��/��=���c9���l���c8B�ϝ�]X�0Z�H�yл*@u/����8�Ʌ�����~ő�POXlq���|Uj�oA��
w�v��˟5�)��K�Qx�O%����aܦ�op�מ���L�,�(!B��.��W2���T�i0����\xB0!�����xŭ�&�����U��?��ِܾY�=`�Zk���Ӆ����[2p����.��W��?�����S8\#C~78�2l�A�� �}���N=Lcߦ�Y�75\��]��!��l�+ZVg����q���t($D�lJ �S�e貓���#5��Υ�pi��A{���I��q�yh�<n�.�����he�8��̻�ATZ㏐�
ր9}�:`|�.�I|b��m[:i��gkE�<Pr�����:3���״Z�Q[�n9:��!,N����	ʐ�Ng�������%+�C8(�G�+��Bb����V���qe��0"Y���a�S0|��U3�۞�j�r��� w^�����`jkdrFt�T��k2rV!�T#{^��H@�ƼY�-�R�W~j���J��7��=>OG�'9�	��j�I���.���������A<C&��!��	��c �
�Fb*�M?]�]��"���]>�O�X9�tۜJ��\�����7t%���yc,u4�9��>����CW#����s��U����0@@p��HA�H6���o$��b��Ƀ���g�2��,�8�;vN��Ce�@��Q����n��� Ox���6�$?�;m*���.ѓ���O��&�T_��<}!~h�`c3ݫ�o9�ړ%�K��ܴB1�e�\=� ��ӂY?�D�墥^�6�.�ê3>�<� �!a����Ѻq׭����{�I¼��S-��j=�fɡ������ �)�g�i �k�؅ЗvZv�C!� "�ޜ1��%�(�4�3��D69�g�"�� g ��F�ӑA`��9��ì�/�*�R�����x �{�"���4���ρKeT�D�P�֦��wZ���C2�%s/2Ҡ���CS���XsYa����F\�lV�\Qn�̌<[j�	��cl��8������@�&����
��	� �XRl�80��z��KO1Y��M\�7�����g4y�����NDH2n��%��l�5�;z:�#����47A�o\l�0�s=�%���9&��p�My��v}�m�����ML�?�C�2��Y"��mW����ͩ4�% W�h�:H�~kָ�P���y|��p8����4��<]qH<�Pޥ��@A�s�C[2Y��XC�@y\T�(lҒ]/�����t�S	���B��X+F�1�����a��	�����0#�Q�\QR�V�Ky�#=�j.��x�z����J�kym��	�����m��=i+g���})�v��\��ueY��2�6݈�=o�6*��ovX�{dU���b��0�R���t<��tf��*E�8���Z!��\CFd�:$��Q,��]y�# �����6Y�[A�}h���Jq|:~^IL.�г�����SF����o�����5���}���o"Z�_y�ڔ�ϊ�)i�&�Y략T�2�sݨ�%y4�Eb�Bp�_�`��'�|6�B&B�͗T ���H~?qܘ��z�@:�V�hΗ�C��E���b5X��I��xZ��Xݹ�^v�����'�����#	�o���7�A5�)�~�������TLBWS29��2s���1�2&�&�:y��{��%q�)��H$['��A�J�3^���+y�}������WHU~���5�մ���^Z�(@]��r���T,���u�u&-a�^;Jf����v[�.K�9l��:'���7�vfKSrZ�_o��	R��������nq�]M1� ����S���c�>.��]r�,�������7�&��TW۵"���ԫ��gi����P��l~���R[nF;����Bg��9��}�{r�{�ܲz١}N��<��f] ���+�~uV���]�����*��m��$̓�>�ް��{��; �Ͻ1TC����9b�[Oq�| fvr���U��H�!��d��e0U#҉���O��6�׹*���"_(�:��ї�TEg�j��XNn��A<���(��*��rM��;J���"֫��U�T��ȁ�S�C��Hҭ��@��3������,�<������Rn�X�{qb�,�{��x��;��O��E>��y��I�;��ƽ��%{8i���mi� �!�R%"0�X�CIW�b��� E�(��*��y#�%�+��F�A]}`K�Lt�V��MJ�����:uY��l�g�i��;�l�|fO����)ُOb�߮��s'?�>�CG�4Ts3W
�O�z��br�,��+���a���N������8�S�U�T4r�ML�:���hKSJ��~�\(�$�g��-���zi�1EܼUۉ]�Yxr,_��g��㹐�̘�Ƚv����k��z�ƅ0f�@�v�:�#��x��Y:A�z�"40�*݈�>�+�����1BǤ4�������L�-e�cD?^�֒��09���Pn�D9l�/|pM8�x]����fp0�5P2�<��\���}��|�8��Vb�B���s����i?����ض�ǫ��qy��b�Z�Dtci>N��ߑg2uo�U��_���� ޿�na����	R~�b�"/y�1[Wz�q��Q�p<7�s��t��dS ҥ�zH�y�g�ӑ���1�z�Ž^e_d�8X%�� ��:�aA�w�jF�4H�v��2�����ɼ�w�M�AdQ���')|���BxaA՟2�h�1ȋsʮAl ���Fe�[����;ɨ��s��zcw��}S���+��d���
'�����t�U6`���!	eif��H����n�+�Q�:	/�w��������j�3���8
Ne!�z���Z'������+��U\{1��ڔ��v���uh:�ť?��U�$�9��0塳*��#r��(�،C�뀢�����8��9�V��{�qq��t��S��<و��K��Gi���YdKi�,�3�q�5�.�������^���!}M&T�A��������_Y��*��n/��/$�˂D��]+q���=L�z�}�};��S��7g�%N��7�(��ӛ��s�@\A��������=ѭ)`�w��f�9D�j���ȵ�Bi8y���_Zc�a���5&0,=�ȑ�RA:��=żK16O����d�7^x������	�wg�K-a����v�7]j_�ʏ,Xg[�y�R�̌���"�*ٿ��p��k&¤�#��Y?V�T�F��\�i����,$�xn�C�˫G��xD$�%��6�������d�hG��b ?�kG��|�K�|0ZlD��]�����t����ede�NY���{�>ƨ5��V�;@�fW>��W��1�0/]�-�tUt8��>�R�A����������`O`��dBd5H�87f<�� e� �*C��0��^�kc��V�p�$3��p�,8h����v��l���!/�IN��jg��*�W�E�Uq�(�w+a��#�.E�?|l{P<k֣h<�\��z����w���-�c�{����$�6�-�3C�N'�E'�>ӗ��I��u�>e�p��`mX����t�N��oSks2:�n��@�"��t��)Uх��t6A��3��5 z@��`^��Ry	I�}h�쪖3�Y{��r�4E��&�tٷ�Əa�vMyl�萭�������խ[����Qb��ϗ��8�O�n��.c�Z{�>��ͦ�D �c���l�:�u�P��\�B�d~�bH<��}K*N��9�?m��$�"V�7o�ċ�:ˠ��0<��N��S<N�����<�E>Pۧ2�̖�Z�@n��\������{S<Lc����c��os��=�����=%k���3���αȨ��d�eW�b�"��*\��E���@͡����;42iNb����{�r
�:����W�T��-�h�̷ Y9FFL
;�H�����AV7��<�R�!�r@�둶��,h��r�饄޿ڡ1��kM���P�G�+�8�Bҥ�˷�Wm�z� ��A�E/9'S��	�t����m=az#$��b'3ޏ/;�� F|�@6�R������f�Р$2Ⲭ|������z��)hY\]1m���i��r��������߁^*)��'�]�+������qi\�(̧�Cċ�!O�va�1���l��=uHD\&;���\m�g��a���
.�*ȄA�?�l���ա���;�����7�'�A�C�D��N�m�*L#�XW_�?�$6Ӝ�e���ÀVϕ�$�e��R�Z��%�t��(��^��+��;��?_a���륢4|{�8S��r/�1��a�*�̝��,�EGŒ���L4V�j�4��*m�S���8�+"�:=R��s�T�T��eq���}}���D]�2S��I�ݫl���}뙰�ٳ�s�\ΌQ�ʝ��EN%���5�O^����4r��R����A�c;��� M�lF�qMI���?$��-������ǫ�έT=G�r>�a*�ձ��hz-J`�8��	�����Ӫ:����0����@���NVH��
�s