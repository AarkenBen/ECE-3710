XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V�5 &�_������\i�AE�.�8^;�"��5�Ĵ����Ŋ��.0p���(�)�^��G�X'���Tx�BKĀ�P�TTb�vJS2\���lH�ιJ�
�G�c�.�YrE�@�Cr�r����?l���X��<�#�|Խ�}a"u�I0?������Ez���Ԡ@����|��!��:pE���.�]4=�S�"l؇|�lNt�ɬ�����g�W�ީR"�v,\	�]OJ�&(j�l�[���y�D�@>�d��1��"۟��0lC+O����[���s�K(��+rv��ą��&^���Yo��jvw9#9ʲ���*D�����c�>?!r��,{֤ˍ�CST�L�\Z~���Z���]>� �#$�Ve��o���ć�F��=އ!�9�]�t�0~�o"�= .vh"��#��t�%���T��x�[�B�9h>�M;��!塅��*�V�tvI� ܼ&Do�=�/�⹟*qPe']��Q\d�b�E7��Rvfm/VO�.�����ԟ~,�-�P�@Q�{=����X�^ޘGSEg�8|K�A�,���+�
���y�w�XݓcR6�w���w&��(�+��-�e���e����n4%^�Oߒi�c{�4x�K[0ޅm�=�1�U��C�8
�7�Z����j3~�sNa�A8-`W���7���p���8}�7���[����suO�ҷ��-g���xyuP��o'�їU�Qh��b0��-�k� ����5�F;��/aR����XlxVHYEB    9732    14d0��Cw&WH�%�K�3 �j�,����i}�W����t��{�������Pp�S�,�ּɟ3�>�OybJ�n�l�p.l7wȹ2}�H/=�M�jq�|a?�Ko��+\FtcS�D�� ��F�H���]��pHy5 �{�0|�􅘹���<�R�0�v�
��9�e��v��̔�[8'g���������n
�؃�����m	a�������:?�P&j�_�2���ygb����q�Ź��(>���i|����o�.T�,����f�n�ѧ]/(��~VM_�1���l�1y��X'��>Cm
���߻���{�K!3�����Q��aO���]����i�\�|^���ө!�ӓi30�M�A
B�ygB��<^��U9|(�c8^V5���]�l=߉��Ԭ�BM��5��#���n��m��Z�'��:���f�����]�F.����۳_�P�'3[G
����q���)��/X��W�K��JvF��"�6��7�Ύ\�l2��q%J��no}�s~�x6�o<�bZ~��_�3
+p�͓�&P�G���;�c��]��Z|��W�>���ԍ��\��B�rui��a��[�N�?����d?Z!���� ER(�@��Q8���r�'{>>�-�qR���	"dįe��m�C��F-6���~�3��8�L�J���������.K�	xo�}q��Ef~�P���hm��w��M1C1�:��e��3%5��V�ĪXd�=IO��i����ST�≼�^<*�\�>�����2]�	V�n�h��Z�$�cGB^�4�wS�i9��c:��$�ot3d�S �L��u�Gd��O2Pu�馵J�������,7��X*����T�� ��P�Q�}��&m����uZDry{]m�m��l�][|7{��E���(���R}���O��M���V����]GA��7��ޱ����q����2~8[�.<�$������E�n�?<�gMN�~B�-��g>���}�8k��As��(f�©��M�(���:EQ[�?֖�	r��m��xb[~���`*SC$\%��Z�3�ATٯ0�o
�[ƞ�p�̴GqF-*���I�yR�/)2@{�z[�Ƃ�hԲs���,�9��fW������2a�|�P}[>G`d{8��4��\�Z4�{�ȫ���jN��HSzI�NQ"��}u5�� �=�0�>,g�S�ı�d��Ĺ��?����w/c�����%C�����7f�R��F�n� o/��	.@wJ�Rt��NV�L#��7x��I	��*lR!����\�BC���T�X/ފ�Ё����9�_������}"꙽~"M�'s/No�;�r����]C��*V�����M�����U��C�k�qp���Qr6Lw*W��oc�peM[�&��9K�:�1	��kn�/S�l��u����M'�m��p��f\vxQ�u�xo��w������c����E��	ۜ�m'�r򰬗��o)L���P[?�J`�5��3o7���Q֝�vwA�[J��΍J���G�)L�WA7�)�B���.{�ܨ�q.(g�A��
Y�dA���^�o�0�aM+�Kd*�N#]��2Q���J�4r�-A:�'�w̭��Ǎ�����>���n'u���'��S�g�Y���#�����?ǲ���`0��V�#ٝVYx�����W����i�=x#��Ԥ�.�����R�ҽN�wAj�p#�Kt��cjNd���Rrg����^	#r�N�q4�Ѧ�`��p�z��ĥQ���D�e��c�b7^�<�n@x�'���.D˺sd���g��2$��z�1]���}#�Zu���s�]+��:P_�&���dtl�b@�%ϲDR*�����%�ux�%\����2������(�ܖ?/�O��.q�pQ����{"�xt���_�T�<tX~�ص&�++w�U��i��k�^d,�>N��7`��=b<r�� {
���R�,��Aa5>�ڛ�^7?s�S�ϋ����2#���Y��0�)�P�v9PH����LG������$��n)�p��+9�<4��?�[��ʼҚ��$�BH�����!�V���|��.jR�ʜPd�� az��"�Y�;c�Hr!����lYT��X%����L�$,��� ۃƴ{�	̽��(�9H�Y�fH��j:ݻ�v�^��	�-�[ᇽƹՔы�	ʓ�ɾ v�g��R�&�}��b��H���(�J���ݱ��Q�
����o�ߜR\�i���ZL���?I�3 L���5���O�V�f�\�"���t��q�d�"��9U��d���V�3�U�j�UB�GPt�ۺ*HJJ�%������(��f/�"�X�$��E�Gq7��C˙��r��T�K�[�Hy�V%�?M�+}-���oI'þr��[�����4��R>��*���t�����\.:]����ѧ��n�4�ˠ�H"ܮ;��@n_�8��S��tVS�e�ZL�Λ/r;E��0����ϫԒW/�z���^7gF�t��G�QR؞p�sq���9H�M��~}��=I,EH�^|�BV�Nz�>�֝;��l�����ZHZS�dw����T�[N�>\.H5.��0��0� P��U�&��g��|�((c�Y�18��8W�hl�K���=y��03�M��LdI�S�7>)j��qiq��_Uf)�tF��� |��8N�;����.��!�.7[7X�.���/-�l����V��'#�Ky���/�P�i���E�Ԟu�v�ͭ�j���qzM���u�zu�A�8)�TN8d��'t�`K�B�X�v1�z�&1���B`w*�Y�Ut;��;�&X�4�|�H�P�L���&z�ٻ�,}���2���R����Q�d����A]Y����tv���J��Bv�stV������0}�ӡ���"��8��2�F蘒���P*�_bщ�ܾ_��Ɇ�*�?���5�)ϡ����1�?W�p��"S_J��<h@���8Zxn���%�-4-�X�2��>�^i��˭E�W6'��w�G������â|����daY>1��;"���B @�~o����C�
e�]���'�<*SFw/@�K�=���J�o;]�j��� WUh��_F萟�eW�mp�(��;q���W��-B�mr\:�*���Z�{��Ճ2]"�ɋP8�=U���9yO�����%c�-�5�c��F���[s����-Α���U6iO��ܪ�4�Vb
�@�{
u	B�v��<j,���ĺ��҃9�;G��r{�����b�{��6o�EU���e�]����yk�V�9?��U��NwG+��@��ڽs�Px�?��t|5�\v��8�ģ�b摣���/�Q��!E+,`(-�r�� i�GI�s>$��\��)�Ӎ�ǌjmKX���Z�}9�sׯ��Lk�~� �Ad�:E�8]�:G��kK舽��W B�4�:��_���l��}�m�b���&�D����T�CBv,?<lᗽ�>�7���壧���y���7e>A��������"�ʕ�����!<���c��>�ˣ'n�i�`����5���T<'d;c5}ړ/å�����&���^�Y�ʹ6�z��%BE/	��L��a�<+'ֶ�]J��ý����|��Ű�-�V��5�!�Z��oQ]�$�V&i�9�OX�=�E�.}`q�=O�H��!6�EN�[�]��#�˪^s�R��,H�c�R��.�(��ڬ�J�QOrM��2Ib}�G����BdAS!%�1���B'�	��#�[���ɏ��䌦�L�aӀ�Q�sb�L`[�\�Q��wJ����L#ơa1X��u�jxAFG�J����5�Qsr�z��T��n*}2����V1�S�@�}��&Y\f�v��"���}�^\�H�����R�s+�{�{C(�pav	���<�nڛ�����ݭ%��G�Լҗ2O���^�?K+X��r�e��NBHR{N#Q0��r}!<D�Ji9����qI��J�5b�n)%����=W�gm�V�&�WƦU� �E�֩���R̕퟽�-Rw�o�/�3�nV�8�6�	F�h%W²C��q�t���~�; ��Ok�DS�X�eL1K5<�}��J����Q�2�,6��&1�g>�g��^s�V����BQ[P���1�>ڄ��ؖ�'ZK������Y�OH9�Go�y�g��z�(e6ji(VT�3 ����0{9�ȹ!�vE+��C`��2�K;��Տ�)^P`X�j�e����^�ph�@��@)M֠P�2��i�;�Q1�QS�;���_�rV���S��4��� �r�`��Ua*��P�yAj
��d$����
��r��K��żwQ���ֱ��ˇI�k�ꢞ2��W�_ix�$���P�f9,`������{.�&�G��ַ�}Z1t���j�!�4G���� Fgݶ�Yen����d�ߒ!Y��&6���k�/��|n�i��:?�.m��"|<��V��ͼM�QE��폇�:�7���C�?`���b�c*|�o��<�i�cK���S(���?��}C���#Y<��0�-����K�h��ؠ�C�!�,A��$00
��UZ�����ڽw���Io&n�R}�\z2@�R��}��Wq��$WN}}(�:@|,V�
�ꥎ�n��yµ/�o�p����=;��Rּ�u��G���~���#i\[^��H �p�_��E$��<��e��\S��Tμ�f֪E�:"v�y����@u���B��2��[;�]7���ڥ��"��ݦ#n��3�b�k��	oc7���]?(�Ը�S����֥���f�r-�X��X缠�;�N���Syn�-�]�2jC�O�e7��>DD3W�If��"**��]4��ń�;'Kf)�9��a�A����%/Z�^�JC7
�;tQ?���O���r�� }&�H���rc���1PZЌ}�a��Ƴ�v���v���~��ȃiЬ����c{d��D��Z��y��ϠوT;�3r�`߽��Q5ۉ(�K���%�����
,�s7���;mAw��
�]ۋ����VB�W���Y]�L�0˹[+'�^K�����{�"���U?[m�9��C;����d�l���"��aO���u�c]W}m��sF�f�Þ$��P~F�+�xC�g�.�N�/#������k,�c9���z��~w�2�X�W���