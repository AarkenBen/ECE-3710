XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k�u�d�/�_n�O���H�T��ߕ�hl��Ս̛��Mӭ�n���[��z�Z[�A.rN| Q�O8��I��!��K����&�A�Q�(�C�.�a�Ƹ+'hF�$ ����x�E]���(���i�۶@�«����@h�f�a%����&$�j�I2&�J�rA����j��u�v ��w�H@�����R���Qd��!i����2N����abLTU��k�S�8�G'N�Q Ʉ>���l"�)U����Y���Q�W�<���#�5}A��h�%������M�\*]'���7�l�t�WI���'����[Ѕ�I�%*6� dŮ�Fk^Dla����*��#�	R��+��)J��ѱ(%����pd��{�f�}����O�?�G��	{O_{oX~m�/7\���j���LT��7�� B�0�h� :[�1��RwSڙ�n�Ɏ��x/N
��Z�¸WS|���Y�O2*�!y��*�J�)��5�
6��T���=�W&��T�!�����^������u�2`L\�W��`�l���sbF)�;!R�r����������;ҿ�g��a�%]��[���n��[)H����Eu��FJ~+ep�B�ɯ��;:�Ĺ�;Y|�N%,MX��;���hypKG���{\�?�F�����n=�e���҂q�J,+f]s�4V�a<�8?��HY���<�1T�摐0^��j=
)R/��4��ߣ}����B���0�K��bҋ�3�%m�h��H��+�2XlxVHYEB    fa00    2480-�;p5k�7���� Y5|hbű�G��wK�f�b������l�jP���<�b��]��%2��d1&p���TG��Y�:����;'!�W�Ze��mX�ᩦ%
鱶SSV;=�"�L�'���N��Pԋ��6�5B���f8�E��Y#�/%���&��zov?�YO�W��F%�L�H��E��؊�[��͖-b��!��R�L��C��P��)Ot�`�O���v�Ti<�o9b�K���@El�l�Q�/�灘=�f�S�7������P_�H�����c�'���ĊF��E�o+�"$��thk��#�"��P명���*m!
�4vL�Q��?�g�b-�w�~�@C��7�8Ȃ���c�'��%�;��}����Ǩ�鋘��P¯w��*:�#�6��I��ᇉ?6H?�#��؆�B������U8E�Yl,S"z?�����:p!hꛍ����2(�X�h�&=oG�T�[�-�@�����Q��+���3���	M�%/�p�S,�*w����υd�&�ьܓ��a���0�a(us}-����\�ڥOK1�� yM�q�;:��m�4��/IR�hIx�z�;�O�-�л��L�7�#P�6�-9�Fֵ��w�NEi׿۩
nTb�'B��������Ћ)���X�s�b�iS��i�#w,/"Q�	���\��kb�o
�l�ۆ,�W�a�DT���wE��~�a��	L[��ۢ4*'9B��Z�c;�]����Ρn9x�xc,�����B��EG=s�!8��{@*k*
T��w��l�RY�Q�0�_5$����R�)^���3�y:zcF�Ne=/�N�`P���ΤA��x� ��T۠�����`<6	����S��yn�A��K���������:��8��F̙�2��5-&S~|�����wQic�]�,rIOJ���?A/w@\��|Ke��U�d����b^ �mdKX}@0Z�*ٶ�G��˜�Z���ڣ^+�p.����R]��W�a��'L�Do���y��Đ �D�-���P~�}�/(�L��8�Hq^i�h��Rӫg� ɏ�.��k�~�sQ�"�疥6���#,a�.����s����J.x��Xx[�ys��oK�?��G���@gX��;�)+3��l��79�<�=	�K_�6} y�W�/q�>����fHb���������-�ǭ�ԓq������
�JTA��vw�l{^f �1i@�W���l^O.�D٨i�6'��^�IaQ�i�x뵲7�}U�e�^��@��p��Yh-b���u7����*������G�h�E&�%�q��vԿ��~����d<�d#����q:�f�g�Y��y[��n����N-]��ovx󍑼)�F۶�0%��
��@F���|��g�i9�(�������\{Z��(��O�:�n��g�5.����c�g?L���	��>z2�a�qJ� ���դض�ND8�^�Śb�����T�<P�p�x�!���`�<�t��5}j&Fi�Z5X�e�幜:�Ӱ>����t�ҳ��h��uD&Be�*#�0��Kp[~x�-��9q+�():��ɩe$N�)�1�B����և��6�w���s3�un����w>T�U���G�jLZ*�[���c54��!Iϧ��hw��2���Iz*��`�|LO`��^� V׋���MN7o(�m[s�����WZ��P�$�(�i�F��&#6Q����r$��7B�bb�K،,����Ϋ6�������-:�۟�*��s��o]d�nEMƋ��d /_VWP>4��h��������A��A<C(�5/������B���;��ţ�����3qЉ[�ڢm����A�H� %��?_�JtkO���z��~8 ��c.3�oA�(q!�ׯ�zi8���N�'W&�E�})��8���~�{����ga�6�e|�l|X_=Ĭ2���(M�|��<%��>>�fk^2mW����*�S�3�릕��A��oa�X��G�ye�T�*��qț�Ɨ�ה_������ү~N���qE��a`5Y�#R��������{~�_��$s!�\�'Ұ/��Y�+�袴<��*����s?��E�vY�CV���2^*��h�s���n�E��u��g�u�_~d�h��9;MF�.%Z�B�~=�F�Le��ث���4�d,>���XU��_���mlw|"�:�%@�q2O_���IM21�˂1{����'s����k�4Hh�tͳi��><�-�8���t���O.�0���0��Qs�C?!����L��/�cnl���a�Đ�-2p�P��2p�l��tm��}X���ȶw�� 1���ⶰ��¯0Ӏ�l�8Ed"���i�^���Ѱb!�; �/k��?�$���aYo�9��>Hzr!��L»��c4�1��]����CE�g���Нַ/b�����gI�0ŷ
��a
�9�8*�F~�vu?��pZ�D��v��q���d����Ao�JU��k_^��bA�X���"W)h��&Rw�b�bP�4<d]Z�	=� 7�ɓ�0`'s�w������GFPq�̙�Nh���2|1�-v^����w��u��ŦJ*?-jH�gR迧U콧MY"Ay=��%j��>=�^We��0-k�eed�_`_iZ_kl�]��O��/¿ꪆ%���M��""+�t2�Ó�[��/@r�T��,���m��t�J%G�g��X���@�&9���	ӧ��t`��At���T@?���D����On�g��Pv�	���!�wƯ?g��<ő�o�����%?WN�{Fhj0`�P�����K�R�q�x<u4h�Pr�J/� �������x;֕I��R5z~� |k+��#lT?5*�?��;5%J;w���sú��-qÑ)˥I�񉰨Ԡ���?�{�/��L�/�9E���̊_'���>w؂��ݷ`OQ�D\nXYm? ���:�mh�ڿ:�ޜ�/?pjS���zk%�����'��F���
�C���������s�d�?���M%��;��[xN���`d�q� �V�V��~�_+�kq�u����z���,*xDf�R�w�F�E���[\B�X_�8�ᕺ�����%vB�J3��T�׼�+d�PK��L9z#����7��Fb�/�:?%RbrXjG����/���j+��:��3���IV"��Ⲽx	w� ߁ei�?���`ְ�e4��O���#ix�ߦDڳQ��y%�A�hVȃ�OD��t��ަ����
/2� 7tfQ�2qѫ{�1�ZCjZ�чAQ�ir
�R���Z�%\�Ͻvl��Fo�7;�v����L	�IC�bq�Zڿ���Q/��h�%�i��ט����!��']�g8,@��K
�C�X܋O��,�R$\C�[yI�Z�y�{1�`�SBU��o�'�wc�B�)*���0~��r��b8V ��,urƇ�J�I�G�#�o-����	oPeϜ���@ ta�[�Xw\X(j#%����#�`��x��ے��nO�6e�iX���zl��2�/n%u�9P���.:aHJCy� xz�������� ����Ec��/��q�����u�����$��|�9��u :2j�]��X{��ӐH�ο�F�M��^���BD1s����(�����L�nIf�h��u��ȇ�|��f���08e$b��V�b��а4q>v�sDn)#��= ����ze0��*�ѥ%�L�E �G��)�����JT�!����4N{)��eJ�d��ȈUޓP��(q�f�/駘
ԉ�L>.���!��$�ǚ}Υ>��C���r�[p*]���[��2S�m��1��{1J�Ө��Lr�O��G]�LӬy��ra�":��H+��f�؁����Y��I��m�[�W�U�]'�X@j~�����W�$k

���]b�����!�>�Hg�@�]Y'�����ՒiJ�Se�K���\����uB�P�{v��s,��c	�Cy
���' ��k�L��(�_�'�-�A~��ei�L������u�`xan�Oa�����wX=�|&<�4+�����S��E}� d8{��Ú���l����y���#*�D�Zp�_�@�F!�;&_ER�����d
$<�m����HL"Vgm|��u�aQŠkT'���k
d�z�r�nQ$8���7��^���`Wl*��tb�Jmk���h�o��Ec��>r�Hf�FU�����ZZ�g�>�H肒���T� ?J�Ҟ��m\��ѡ/E �jHxx�a%����|55�3�d
��J��?�o)�:����i=td��j����K�bYy��l%S?�h�e@)
��L�x�:BǷ�/����Q�zOc(!������@M��[mJ뙣*B{e%®(7��t�Y!R����`߬ẞ�Qy����.p��'���wAJ/˺4
�<%�X%kn���:�X�z��;s ;�/��x�:ر����L���a���HcON]Bb���О�GG% ��	�N�t=U
�2	�/|ꏼ�\�#�_"�W'Y!%��Iuw�	�u�������v+�������J]�d�]����'?8��l��9�ʵ�F�-Ϳ;�,��K�rC]��79X#׍��aS
����,N�"����[
��E\�h�J)�T��������ٜ��>q�)ɒ�Զ�]d���*��^��FR����!S3�_��)x���T�L�j��>��\Fw���������k����	pOj��<���v�Q�d�
�Ͽ�"��QjR�s��h3�-��P}� �����`x���[i>di1��t�v*� c�7������EZ>�������X�ԟxZ�����7��Y5����t�?��h7���b|s�8I�;�n��wN��`���Ṕ�ķb�� �te��U�{]���7����� �|N�A{��"�P<�$��p!ُNt~ţ�6\QN86�����U�A+�����f�hO}mr�A��؞ۥ��Jl��)FYi�����-��_�.��!a.�#�8�V?��➥;Jq�1�k(�1�������>�%�����.��_����5cf���on_,7���/l�v��E<qA2�J��wt�"�qo�T��G�v/4��'}[�Fa��9�MH�ed����i�إ �� ��nt��4��(���UNZR��O�}*r�[kB���i|��-F�b*u�������ix�*�9�r��xauz�0,�g�!�+ўq#�ՠR��ll���x��&�pԀ���~�Z��BL?���#K���zi�eC/գ�*R��6�9΍K<��֧9�wd�'�&�~d����xOYl�ކ�n?�c]>���-��l7������Zok��Z��a��˝��ے������Cы�ZpK�^�/צ���/�d�8ɏ�q�I[�+�Ǐ/�h7V�-��ۑ�^c�<�n��C���Y��,!��#� ^�C��m���U.m堌�~`7`�չj���[T҇�*\}�����C��sId��W6�u~�FP䥫\Y����K�l9����Rw�Ι�/9��9���@��j��KP�tRM�?�`j��=9�S�b1�P`�|3D>S��Rr�R�FU��i�����yK��PP�U�(������;[�G���1G���\�^�m���&�Ji��:R�Aha�'6�( �v�ޞ�&|�}�rz���Rw����i��n�%n�m��/I"�9"�7�y��~ B�I�®\��r����'�F=� 猀Sp/�jK�ܹb}��j��$Gl��i��
'��r�4����z��4��t����#�#<ڗ��GWz!_t��*/���4F���ԧ��?OX�!�tD9O;�%FN��'"��B���)K��[�)SEz=mj�y2+�&����ҁa�AP�
��6<�#/#H�m��G���5Z&�H��":*.��W�W�փ�Ȝ₸ӪJ�Q�ĿiR�g���{W��h��_m��R��b�ku�`W�qO��x�F��8L+���lU~[V�v`�p��K��(�4k��o��Xf_P�����������3��1a�/l����ӛ�!�_q?f�����Ϳ$�!o�c}M���̲}�2�V��m1�^�jA�m|���o�2�y�bȞG�'-xt*�G�� Qم
�_TG����FXW��
	\a���0��_����kl�7E(��o���zbhF|��Wa�g����m�18ֽawϑiݶ�<�2�w(?-� P�?$���d0�A6�C�Ǡo�g��LD��{ݧ���[ ���P�$e@��N���	�;'��F�Z�ex�����׍���G�k�*��P��+�0�r��2������yA�+����J���(��r�R\�?�D�ӑ�:V��4��[ˁd�sw
�qbT��y�7e�p��01����;���s��H���Yz���G���� ��[d��w�^�(���/v�ќ����'���Bǌ~�+ߢ.��]!�y��֊s+P��ݛ T���B椊�eu�Y3�kBV�=h��=���J=q��reݭ
u�Һ�I-�C�S��t+���s�p���������[3d��_@�kƒ�� t��5�a�R� ���p@O�8
H��4w
��B?'L��-�_�*��Ba��T�
	nRe�G�d� .
L�������	h��4�Ne��k���������=3�<������Kv<y��+Id�>g4 Y�����1����$X�����eWkg6��:'� o���r�i�-�伓�yv+:�apw�<�-�E�Cj��3�����M,�GV��I��
��x�n:,+9�:�*6�����W~Ѭ�J�A�zH�����v$P*���#Ik�|B7َ��lk�."�����yi�BVkx�y[T��-�%�z,�B*C��>��:ߗ-���$f뫡���g�q'����/r0v�R*MF���u�p��
1$�����)��������	A]��-x��)Es�l��
����n��T���^2mtu�j���v�"/H8�L���������~()�@щ�G~7���C��2��6�����v~7k=���P�Չ��u]W��K)���y:l��Y(���)�l���zB�C@SP��P�`��������|M-��m���XCA�S�p\���/*�Ή_�� %fGl��1T�%���?�:v���+��͗Ph�J�	U���u�{�c2-��^�_���NlK+p1��d�A�o�hp0�=6��F�
GT@��9���o�յB=�uI����ݨ��\M������0MDF�#Ӥ���xbwd���~yCzȨ���X���\����
�ڋ���pʮkGD�"��G������)�4_�%��m�0� p�c��׆E�fWF�ԍ@ˮ4�nL_��d���pu��V��ֹ��S��ok��В�c B�l�K�������nEE?R��	����R��QxEnE /	�]�QhqEUxsΊx�t�["�����*�-�T�<���d�ߑ�p�W�c����W˺�<���\0�q�����D�a�%��w?�dm+����Y+Mʸ��a��{�W��:�y��O���=�W:�Ū{�´$��n-W㯯��v%�As� }l�jLV��w��\�Xr�&���+Y��"+�
��V��O���u��{AM'�����s&�>�sBx��(���p@?J�������oF���mm2����\�O9�M� e��K�J~����""Bұ���+cƖ�]ym1p��g3U�ʌώ�**���T��+���9�0��@x�<��;���s�JȮ��ѓ��< �$�/DKr�+�~��u%X�,+}��f�@0 ����쎸��0I�zP~+�ɭmyݞRuP�[����F��R�'�6Ll=(݅��m�;)��؎Ϝ[�A�z���_�&�c��V9]st�n����4��X��\�tv����z_c����g��R�ѴC CUs�z���K��p�`�M鴇rB���>|���d�p4� 
[��
��C�d{�UnZ>B��kk���ш3�q&$��Z��vX�y�.k�c��!���ڽ(~�R-b��w�ˌ�ip��]�#��V�sL�+���]j����l�w�dG����ͳ��s�3Y$U��.B��D�f����u�JMA�0@d�#0�����w�6������$�Z�ō�G�}J��>�i�F��/VXX�����/��d�'�R��=C{�>�7ۊ�0Z��!�O��QP.���A7�R�mT����1��#� ��[� s�\�����P�c8}@�yv���JU%�iS��ɿȭ�t��q�@g�{#���-��S%$P�$��,s$�1 ڀo(�>�MT��ɽ�GO�Y��0�L��O����I����J��.V:b[�a�nԩ�2)^ƭ`�f?;��r����R�^�ݍ4%�c���Qr��W
�>Dy������[vAH�.k�Y�︃�QՊ�ӑ_~��	�a���4n�]gA�ܛ���%��A��8�}m�RA��o`������3�(�
6��"l�����C���;w���`]��)��I5�B�d���}�J�3��g/�5��1���g�������x���F뇽����~yY 樮��W����<jB�lO����u�G�bnu,U����i�
��h�?ҷ�J*#</*mh���#�f��zn��������	�tm`�7��6F�<��8�J�j0����j���S�����\�л�2��� C3�(û�Q�s��γ�+X B����L������j�6�[�z�y{I�]���qi�)�s_hh�A��ar��dI�d[��3r�����J����I06��_������Z�\��h�'����M�D6�<θ,.��B�-l?'�$ﭠ\��.l��BȨ�A/��u���Q*dPR��p��h���]NHf���`.m��C|�=� 1zq]�A����s+_Y��eI[�F��$�"O�_��_U��H2����	��w�N�+͓�I,��K����^��Q���P�D��.��\�,����s��}�߹G	|�MSՇh�����l�qIk�j}�J��X`XlxVHYEB    964e    1150��Pp��|��e߉>Me}@wk�vز��%�$��~����*��U�Z_mu
��m�"6��������|U)���z�V���@H��x`�"��W�i�a��3��t-e;���Ҡ�bTO��Պ8���'h���cZ��.
ޤ!V��!��(��"^~�����g߶�i�����7 ����CÞ��3O�������]�o�����@n��KcT�Kk���ֲp�[�&�m���S���/�YU>�5�'�Q��������S�+9�f f�����F�(���@��|�GC���f(���qf�v�ΦV��;`Sc�)%0#ȕ����VI����Ia��f���;qZ`�Q�3�����@;^a�1]&��:�L{ݏ������Un����`���#�TzP5��~2��c�����������h�/��yޅǏ�� ?5]�u[|���LgJh/�������
��8i^�>_�~�vJ���O�'�i������� ���a�A���>�_��
�]Hm cN_��<nU�q�>����<2�.!�y��u�x�2r&7/Pk���hq,�noqoË���-�n�Br�h�O��a0K6���щf���+Ą�'�+2ts�JZ�d���A&��~թ�HV1�A��&���|J[EL��)-��řֱ�1����ND%�.B��{	-C���(~k���)/�aAqb��}�S��=}��Ӗ���K�YW2W��l�۰Q/1�iK��vx����V�U�c�Y��ՙ5^hݓj���T{�ƒˑ��(�Po{��Lڜ�*0Z4Џ<�&9M�낯~��l�ڪ�$� ��j�sc�$$���"�'JN�w��Z����Y�}iP%�����(5`�R�Un�>���8��dI�t�ZRLL�sg��B�͝��m0jkuչ_�J�i�Ac��1�ڟ=5�H��	���е��_�f<i}�@(�2�5�o�r��d���T"�a�a���VV���p������Ym�$rϛy]�	� �zchc�#X���[�OD��y{>�3lK$P��6��y� �25�a֔�c%�dJI�V�p��0�w��o�밃��}LǼb�ņ��,���z���@y��˒/�q# 0N\��@�1HK��@�|H&;X��]��7R���ـ�m�MX6�����O�m$߈�X���~j�TK"3!%X�UPn��ߙD�f=������P�4r"���(�[n��A``�A�����c��s�{�u?`��o厙(X�
����q�Ӱ.7YFu�˶�%�&_��󜽹��Ƭ�ZF��:N��-�u8]�lm.�o�fP5��[-�_0(��ڛ�,��D�n3���̍	/�o��k�tSj��;!,��:Y�@W>��g���gN[S.p9��vU}�t'co2�J��o:X�s��$���3	�����t���i��52=M{9q��[}`��HTF�h�ˁf$RM|�y7OCR���
�g`2�����.��"5,v�_Rˈ/�����K�BSZ��#p�����?�l�0,��\- !�"�	RkIy�򹑛������9�}�`�V6?2("�tJ��D�`p��i�&�B?��3C�˟Ԍ�TUd�e�x*OH �K
j��P������w��ԓKt�	�1BՎj��A�2�7�z#>���	`�"z^�<D��p�r3�K�@�RV����+�]ֆ`v���a�!d%�i�xH;�]��чb����7Wj�L���2�2y*�Y�x&��mq��=L���S�5�z_:p�7�cϝ�'�������-���B�G�;R[�؃ꦶ��"E�~�V�G]����G�Т�s�C�/��A��*� �@yT!�w��} .����j/̒@�9t�]R'�.糱4)�mE��lͧ�Z�ͪ^���'�ﷆZ`��ҕ���YҜJgyO: '"�S�;1���j�a5i�x=Phe���M��11���=�M�{x�����T˚3�u��&�	��&nߞ��PA�?�}SC�T_���+��IH�=MZL4�d�b�K��(���~�2I�Y.��;�0�T��s��E���p�r�6�C��K{hU��x;��rs���B�¢���D�S#�_c����;���
|[.�=��S-Ϗ�'�7B���I�Ȇ��]��;_��0���ݸ�+18Cɛ3�XkEHx�h�^���&?\C��S���ꥌ�p��Wx�%���ܛ']+T�R6gI*��z��?׊��c$X��#\|�hÈ�#c�5����X��.��/c1�y(�����akĵ��4��RC�{fJ ��[�E:���e3�vׄM%��o[w�f--��rP6v�zjo�F~���xڪ-?�<�sh����^
�?!� �8�*L�@��*��%b�z��RI�mӥ�Jc<?�=�Y�d7*i�V�#��:�0}rX)K%M�3D�+�`Zn:�b�	p�S�șb�7�|��5d|�'{'�̲l�G̍��^����i���[e��B&1&����S`�.|�di���ղ�f�98*]~��W��@@���|'�z�h_ms	Xط>�˪%����
���֚I��ҹ��>x�Y�)�V�{L�l� ���o�is��@��({��F����"+�}�DLС��Nb�4��ݵpS�v"9M��;��P�DE��P,�*���INpE�T��0�㮬y��z�cP�@
n���ǈ�!Ie�׸�2ree�ċ���A�3#t�k��C�P݌�U:�;.��`��H������̺�ޜ��{Ep�#$����E0��"$�,[�_���Xka������g����R� �>f����q,�SD�nQ��9i�iC6��F�I��Ę1�E�]k�Hp}Hn/\D��f�=C��z(��J����n�
9ΐ�}�T�E>�y�A�3kRS:9�z#_�f�X����%�Sj���q0^D���~�x7d��H�kĶ��T����/$|��޽�,�Ϝe�@�'�!�բ�e��}P4�Elak���.���HZ��nԎ[q�?�m�!��{�1�|v���r�!�n�����ȵ�ʨ��ʌT=f�#g����AO�=rѰo��A�H�8�^z�U�xˋH����l�͐g&X��# �`�P=}iEy��4�Q���]fS"��X���+�T	��Q��֓�Q���(�i��v�)pܲ�j�__���_S쩴"��@a�F��S��s���mBn�eT!
�^sWT"F�'���Zʸ�˿)�ަr�4*~1�r:�!I66$s�r1e(ZdK���
i󬱥I��GZ�l¢�t�G/R���<z�컩��Y
�ą����h��vtk}߯ͥy�ˡ�JFr���=7u��g�e@�Qցlj
��P�wWUS��T=yq\���r����	�'eH!�3Jij�2�hԸ{�/)<��E�@r��tq���
܋[5�zD�_�P����]��fŏ�-�]�H�1�w���>E�����K0;U
���c��`�
�;f�MlEI+T�,7 �ߪ`*�n�/LG-C�H���b�O�FE����۴1��g@xR4
ԁ�I��Ο��\����eP`���R�I��#��p�ӄ��Q����3�[<�-�zެ_̿a 1���~η�cR0��?XyPM ��x�6��99~ֶ%a����9�&x������P��{D��W5�NL�ǝp;�P;x�,���cjB�BM*T�ClH�j׊�2�dE??��=�L�D�ٗ����V���g`ƿ���,��[��S��J����"��MeM����)�ַ��i��qǼ�Yp2�a�9B^�:��R,�T%�؉���N�-� ��d�:?��pK�������	c�� /���7'��D�^����RD�&?~1�f��]/_�CC���m=�e��R��m������v�^��t"��:_�ͪHx��}�qi|��o}��_m��%��^���{��V�߰��p8\�D����)�?
�����;O���d2��Ս��P�C����vw�U�Mu��k�9`. �gB�s���]7�kY���rj닩�V'"�BM�Z-5���e\!�����W���S�����K��d��p����&[����C��M�Ja�~�^ll��j�r#��z�N�/�x��&����/�Pn���!�[v؋��	��>.z�R��9�֔dӈs�P#�c*�Ѷ@� ����hH.�L�l��+)�aǮ�gye}�¾�x>��;ZyD�e [�0���B=Oʠ֝ݠ)W�b�d��c0���g��X�p0�8�ѩ��7�%���o�
�Vü$���j?dB�OiEߊ�ƿ	�h|~3��f|�"����+3o�����*J.�$�����T