XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������������ll��y��vՃ�t�J��RHλ>�\~��s�Ey���Il�IϬ�IP��h��Ri&O����}uhh��9e��$����S1�X�NcL}�T��'��;��Z�#$m<���y{�4�Sw c�q���f�I�f�>����Z� �9^��t7�GT�jB�%��@ʀH 究\8CE[��x�iR�BB�4 �sJ��N���1��O��<c��+�6,>��F糋��p���@x�X� NݵB�����S)�3y�Df��Q�����QA����NH{j��?���%�G�L��2h�oc?t��T(\����u�-y)];��nzV!���66��%�[ �Ԍ��g��j|]��`�}�_?2��.�g��rzH��v���wo'�"��r�z��緈�P 6"��ibu3,��*k�3W  �:��P���A��;7U^�c���-�Mk�����W�u��e�좟Gh�g�S�H��9mc�[t��
8��ӣ��:�]��靯E����v�k����}x�cep�?���bV�%}����L�*�n���Pt���u��<�fNr.�G����S�����g#��3�Oh��}�ez���)r1��"݂3���UC&	�b��-��̒�;'���ra��?Mc�ŀa�@���N��%П~S_���,�����+ZgM��1h�\����ߢ���cad�}�:�ihib��l��O�rϡi˭�|�1�W� (~{ �<F��%b"nB"?��XlxVHYEB    fa00    28c0��No��.��Z�k5�Y���q�� ��kYۆ�_��V�k��I�����߲��~0�:�R%)N��:F�c4tꟉ��W�:H���p)s�|]�2fP�&���B�!lWna�]�~³-�(��D�A0�#���W�56S_�3����cܴ\�a:��x���M=������K(�h�4~�-��͑c��H�Z�S�w�v�h��iԊ!���Cp,&�����o�k�8Q�q���Κ�8�MK�^6h	נ��"
+1���7;Sqq([���z�Z)7�K6,lca��NH�|t%�)q�z%���fmMq�g��-`�kvZ��w*<�gM�ɿ�N�8�8 6p�����[�Ps����g|S�c�8��y �E>�Y�
��f���xB��r�U��z�d����v�b@�h��s��A���tF#Ӭ(i��×��nȄ#{68M���Q�떦Ӆ�ΦcN��U�	/9�Ou�:)�s���B�m.tgAA��rA������C�m�:�l����ue�Oo�6�����/U�'���d[%�w,��'�d4W��A�lu͌��BD���=����댏	�bEAB����X�{U�1��q[Οȵ}�6�et�(�^|��㕜Ϊ��Эua��nK��0d6y$q;��P6�ɖ�^��!:n��ICA��7���ո�t5�5�R봊�6�<�;RҠ#�J��+uq�����VE99zm��;�C��.3�ؤ�$�NB#�����c��]��a_��u����O��ǒ1�}(�jr�8pn[��6�J�:�0t�"cn�����=֟ؽ��]{F2�=����om��w��)?���Z!��yc���Bpc���	!vczf�rB�'�HM�L0m�~Ț*���1�0��Y?1����cw��m���6�V�#���W�y�-�0���X+���$/m�=�P4'4[:�|ڻ��C��C��x��'����_���W^���zy�`�w��}Ҵ��:�)�������	Y`^O�/����}��K��� �=���X+�!w�eQ�>x:���71�s���ޢB�V��;�7��?4`fVDs6%@ �?���(�?,�X��>W�~Q�0�����M]F$ēY�)��"��)(�D\�¹���Ǣ�񡡫�\���ԣ��{��ީm�U`��p9{�ޭ���RD�Rz	��L�XeV�)��(�IvUƩ?���m�D�=y�q�S��u�X�in�J�]H�x���y�g��O>���PH8�}�p�������2~@H }�Jy2|s,�4ܖ�VSF�R����["�v�^��\�a��|ǐ���luӃ�����#�d���1���}`��j�l13U��+���H?B���$��K�+�z�L7VrPe���ؼv�9�?a��_r��3���5K{����O�)�D0H����2�/�J�d���G������0jO}���81��L\ҁHI~���-X�`d��l,eO�OɈ4Q>��;ʸ�C�
Aι�8V����i��0��0���6��`;�ǆ����@s�C)�M��	`����W���]t���]��ξP�`��8�W�<�&�Bl9�z���\��e|�I��A���;��Q�*�c�m�m��ߛ�40�`��ZȾ������nS5���-�����R뜝��+]�@D�K��i��ێ�(���G���?堄��k�n��)*؉X�p���^Ab�Z�{�4�L7)�C�}�+Ji���J�kм~���:z�@b�8"� ����lg�<�~�Rp�]TW?�9�k������6�g���(��NQi�2�k��Y/�2����:v��ڀq
�p%�5ӊp�f���t�
��v,O���=�J@�SOX#�;J�d� ˮ��� �s+�b�:��X�ł� _��Ƌ9��b��OQF�ŕ�ܵy�P8P��t��Θ�:W�Th�A��� y�d��>��{2^W۞=8��)5}�����Ğ�qy�`-*7�ʷ��Y+K�� �_���v#&E�0�A�����C�j�V�d�����tc�$��*]�c^�̀��JiY��E(c�d�s쮯����5���Ο:۵㘁��li�"��<�v31��p��R��@�\����%׵'T�!)���f&s�c�3M�Y7�v���S�f�{��u[+_��}�cq������z��,�k*TJ'��W�8��38�@bl(O�u�>�e��&�:2��D�"���k �̍���nc��U�OMў����R����24ܮ�X�y����t����Y˛�.����Gw�B*�N����2�̲��;���+һ����-e\�-ê�^d}.���s�����_����h��D�A27$�*�J\�b]}��h�c�������A�˚�4���=G�=�5"���D@�S������)x��go#�J�RkTκ;�Xǻ��B`�4���ǩ������%�^��5�ݙ��g��kgL~�e��	ŷ��3�
�i�h��K	�s�.���<�����UD�&?k����= ^,vV�?r���]��im�1@>$W."Կ�ޖ�0��Pd$�t`:����r�2i���т�/��}���9��d����٫��&|�?]�'���T���D�� ���_([t���X��ڜ��P�أ3��g��X��]ѐN?�΂�{��ʙ��Sh-��®a$'ؚ��+��Sy��̩����&b���ED������>��1���o����#�����݅z�Ȝ^�U4f�)@�[���v��jTǰ�$sY��VYJ���׀�,�A��,ǚLZ.&����N, ͕�"���Wԃħd	؂�_���r�*ʏOdF���s�z^F�I���~& d��/�ZdO^�aq�^�À���}4�L�ߗ�kЪ�>�hbg��5�u���66�p��oAxU��x��Q�r��+I�=8H�����H����R���(P�˒�΃h�y��d�c�T@�얿����]�QN��//"������Y�ˌ֌x���?��JƂ���釋ˈ�9��]d�Fx؝�H���Ä��!V���vB�~��Ś�&�oG9��v]�-�-T��(ݟ��i��T�[�����Tv�JC������`����@�2��h�+����S U�?R	���b�b)�PCЌ�Sd��03s��ƽn�RϬǻ�ׄ�ŧ�+�.������[�s�����b�r�����@��.Z����=���yH��2�8��f%�.	%����O�e}�/�xZ���w��ya�Т�Ԃ ,��H���c���O1�L4��)ފNa��͟|W���F�z���C����fD��!uh��5��G��6��]��CoVg�����6�J�Q�I/�Ifc��,�y4��z�X鶣�)I)$ؠ�ZI��g�-]�Y��`z��D+�S���R�`�cPĨzK�$��o3&�0}��bPY�d��~��*J����9R��6p�Eyk����&�l�_�� Cbc����#�vh�;��"ݶ!���k&�9���!Q�X�	8q]z�8���CPv��R���A�_I����X�۳ie�:�I���G]�@�����Lh���)p��e6��M�7,C��g��x0�ć��	�1ۛ��1.��иS����qi�>F�j=��MQ�{��A�l�Rٔ%�'��{��-��8�$����<w���j>}��P�XI��FPND���,ꆟ_���܋Dk�)E��d|yc��UN�;�lu[.2r�����������Y^>��׻�[�=ɾ)�R������R�u��i0YH�2s��BjK�\\f�7MO�T�d�i��(�@S���C���	�މ�v����V� E�Ke	�B�C�ԈxN��:tޥ�+,�$_)oH��=$O����?��� ��v��;%�y��B]���4�T�=�緙��s��I���z?�;����ܬ��c���9�Q}����g��V�s�Ҕ����^H!V�8h�_:1�Ά�X�����ܧ�uk �깳�JIk�)���l.�uY�4����|!�I����j�d��bv�������TeV���N�l_���vڏ�?o���yK�R��\M����t詊��8�?q�e?���fxg��ŏ�X��<�LyU�Q�����*���h2>)�u�q�TWgzڻ��b��#�i� ���
[5�',�ϖ��6����-�O����3������H�:��(��),�������m/m�}�M�]?���i��m���U�>m��, ���]"�pZe#�����RS�2`��t8����c��*�k����k���0�I����+fl��U^����D@�;fJp�y��5�9�
�����:�h?=�r�|ov�����æ���gjt�r֫��!k��~�B��܍ߨeC��a���x9P'��	o+~���x�
��j�����C�`�8���$_�H
�p+=��C�t|�\�p=kS����	=�y���`�S��\��0tp-9�YE�a6[mx�	��R���xC�*Rl���}��o♀�)��U��M�HI�����"�!��@KF1P��E
�����Q�=f���@���J�Ɗ��X�m�aWNP�Q�8_oW�Q����BiC�zҔ��IPd�%�f���4;��xL�����̎�h�m�{A�ld���.���D��$�� �,Tf���֕�CLZT=S�\�+.k�nt��{|�ų}cݓE���i�wK�d��z<蠘>����RپS˛�p�d�ϩ�zoJ�,ʫ1{z�S�m8��k�v�q�AV�7_h���L`��&[�*]���ټ'��!�z�(������5A�C�uC�����$ �'"܁������"�킙��n��<ր��L�&G�F�]PR`��GmD��u���Ό��(� �Ca��!.4M��G�U�PP1H�p�RF��`��E�M�r>U�ЗV��r �ٌ������?^����Q=�b=�hO+��b�t���+�r�iwPj�^�ـa���wv�EFڻC�M� 
Zi�u�h�׫Uʔ��u���s%�I 1vyo��%��}7&B����}/�EFd���uS��y@��*�������[I�����3���׊���,DX��ZǬ򼯿3:���E8{�-�i�jw���	��;7t������_# ������e&��<�Y�e<�wq83�ͨw9�P"�I�x�f34�C�	�{x�O��mA��F����"G�i�"�x��4�2����p2��^~���,�\�btJj�6����g,�3����;?v]9;z��#���!��I��w�"I������}E)�BY��/R���P�����)X5=!߆1�s)?���H��i��m���?'�⤓\�3�䙒�*��[[��A��
��l+�6NͽPY%1n����������-]�v!Nt~���؉����!f@OO�� ���GM>�̢�J�,�j��Ճ��!0d�ǧu�o ����^U�1�J�p�d�6�M�}RO�_�oIY\\���w�0�-��{�yF�a��x�,k(7]P7��|b`|N�0�����x���d�JM�Z��w0�[߲�� Ĵ�$��K�sl�lUp��Bo����lD�����\=?N�d���=�S�T4�:�J��KC؟]}O���F�*L��0P ���H9��R=T)�L5��S��U�Ս��E2�%5t��]�����*_��]�>{��AY��8H,"���'7T��k\���<~��g��N#��z�h�h��6\H��q������y�޵>]�YY�oT:9�$�Q�|�o�k�IY䃘"�Bup�q�/���J֨���O��S�\ڮ�������e��	Em�/���}_�z�'�����l��c�\z���Jٹ��(�.t{��"�_�ҿ�h����֖��F���O2>����=��V��Sv������V������������;�T��T�����?�܍tG���t�)�"�^�ɘH����(�l-@�QZjSt���9:�K�e싰8t������@�U����	y>�Ռ'��0;WN�g �maN��ob�)���5dmʢ��R��b��9W;��ӞV��t$�+ ­_-��j);����_�lzH�1� �\�t���2?ǚK�ٮĽu
�Y���U�!#���T2p�z�l�2d]P��+�|������S��z�>�'��K	diˈ}�q��(���[�۹B���JX��_��J|��c���UD�1��V(�/�9@_�Ro �Ŵ+���Q���ka+6ELޞ��jX�I�X�oq~�ٱ7�.�)��,o?4~22P�
��������6Ba%'�iȦLn��t�Z�����oFm��+v{ͦ݊^P�P�m6��n�����&t��-���uq͹q����Т��������d���Ƹ7{����9�6���b�$ԗ���2ޯ���;h���bJO��w���ꆻ^@	'�u�e�v�z=��V[���&�;PE/DXW��oʝIV�)ZS���,;.�}��N�bʩ������6>�R�yZ�{O�B �Ht����\z&�P1A��6�ڧ9�z�U�E�!i@c�����x*^5�ԧL3�%���:�xp�����ȉ�L�����Zr����"���}a�.}JR~d��b�x)��5}�H=_<΀��F��2vAz�
�>��|ԾGY����9�(P�:���1�E)�����Mڈ"����ml[��a�?�J��4y�J�Y!K_���L�Vjޜ�&Ƞ7��Z�4y�ܗ��i ��BT��V1i������$`>vô��-�n��X;�08veR�T�&Y΋|���.ɰ5�qL�o��a���&><c�0�ƥ� [���p�"8��B�-i�WM��.e���zf"���6I��څȜ���
\�"��
�Gf/w6�z�U���*�Xi�N��F5PV%#���,1�����b�#כ/��)fK�]ɲIr�.T�qӽ�[dN�v�lw��?�Q~�)"�x'ވ�@���۴����W��h.��>t�}mm��)����t�B�7�xtns��D�s�z�����n9��\FG��	�o�s�[��EV�t��m���7�`yXi��3Fp�0��0#3�ȣKD��j"�|�]�G�HA'�1�T.�t��v��Jbm1��C�ii�'ՕfҘG�w=�zϨG�p$�+�
��I&Mf��o%@"\��3`�M�k����b\nX�lm̐�X�W҃G��_�/��Wgp/r<�՞PV�x�玈t
�^jI��'��P�����2}Zu�(�sG3��UVf�z��˾Gnh���V��RE�5���Q�}!�%��}�Lr���:Z�����A�Y��#"�hl������-�(}wx�2r��\�%�k� ���,����t��
x�L���!���]p���d���QH����Z�KQ!6���6=-�~:�#ū�Lm�N� �H*#��J(��h\��~�eP���j{
��L>�5`��G|2���Y��`'3�k墙�uSH9 B럟X�:4����~p��ʇ�q�F�[kYUE�k����>KZ�\_��-Sɕ<ݱ�����{�bJ���w2,��:J�5���<��H�X���1�;t%�~8����O���R*�?�7�D0@"���eW��Y�����'(�:
�!�7����G.����(�| ��� �e��TWr��t�cz�5?�g���$�DCy�NL�����灠�=x�Y(��$4�έ(��jh��|y����J�9�hfNC�#��	��P����)0h��t�]��Q��Օ��ݚ9�t����-������
r�B
dO������(U��R9/[~���>g�@��Zʩ�̚�ofD|W�Y4*.f�
uTͭR"��̊�[u�f���*ͯ�j�������i�8T�
rkS��~5<����G��v ����lB�A�1�n�ޤb�ōe�q>���R�M�zu�i��%��a�Ej��ڋ0؂��G�1�Wʞ�v3�����)�'�%��ȴs��̮����<�m�5A�A��飯��~m�l��X5��,$0�f4?�hð�]��݀~��+�Irg�Q6nJ��^~��I�RL�͓2*��;P���eN��k��s^
�hR!<���L��0[xN�h��Jӽ�~�^��¿cU�d,Ж�Xβh��ڔ
n��*���B��=��y?ů�uw=�t6�<8s`�g���wO�j�E�=��N+�ۧEI#�%K��t�����>���r�GQ}:�VX�oVn�b���^A]Ԑ�?��lw��C���tA����<R��p?[t�z��$F���e5��=�=�m�B� �����*�mO�/K����1�y���V&����ýdv�O}.�s���<�⿍G��x���w�	6�s=P��I���G%��.w�Ž4�٪gN]]ʂ�UO�!ާ�!��֗��'��O����j݀%/�'��2��ITsty {�w���x��!vtG���'���Y�KB�=��"��xd�M�ʮ)\�����odv��E0��I�L��B'%6��G��������V�6>Y�N/��#4<���˒�X0�Mhg���J"l��Q���4���_�J�*	��͠�:���1�{���}�Z��f |?�@C
\���8��_6���ѧb\c�>�5-�È!�^C���iBEE�b'2;qzM���&�$KeC�E%���>v�d�`�)�c���d7��X��Sy�g˻�g+�FpO/w�0��lt���A_�x����Y������p�3
S|9�׆%��<����ѐ�Wu��{e4����1g�k��Y�t�H�1�����9�j��r�!*��B��;�S�Vsl .2��gz�ȗ�9-5��1�\s���d�o�6����2V���J�V/[��"6�	f6��7b��m����t�=�5��]����+#��yЀ�f��d m��&���W	xB7%8����Xv�#C��L\�a�.�2��w֧ǘ�pq� /d:�ʠ�lP�4٠gu��Vy�O�!�U#��
%P��0|��c[,�h���K��ٚ�ܻuO���\v5iEެ{o64���$���9�@����O�����([�&��K�ٵ�0�u�Y1b�u�Wy�|����M1�!�8T�� ����O�W��a0�Z��v�t�a��8c$O�W�H]F�9�s�C�!)]�.�2�>�Ȏ�7�[�q�OK0ǖ�g�hA4/Q��"!6w�~��y�&�E^͉�l��>�ځb�2�I?��N�u�������_*ҽ
��?ݿH�w���"b��wR���P3x�Dap�w?�mq��ԡ=�-�Zz�S�/n�0��t���FL��5{�2�F����q���O���t/��h�'��)�������I��ަ��sjg`��3��_��6����TO��@#��|��~2�bV�t�d2��S��4Lݲ#��۠m���*�@<����!f{�!�I|�� �YSgix���M�@�Wc���t�S�p_���q2�W;�?n��ػ��R���ɘ�)�t�"?u� �S�z'jr���v45>�7`j,�Ge+|�]G�������8!�X(�D��nJ�%(�1��И��J�J�ROq�X	mTf��v���#*?Xst��,@uF$.�-������Q�����_���<`���ٰ�z
�d�m�GUe�a��a��LX�;�r,8�/sfq�0#)�8'���|�h�]��jc�(z+�w`�z�4�*S��&�H��L��.����ٷ,����DE�V�_��>K��F��E����y�Z\>6��z	"���)u�D���z�1{sĖ,��4�O�D�F`�J#%�Ou�����S�s4߯��D�p����+_��Ŋ�E���z6��x����Q��;��9�K�=�������m�G}��DD�'P=ٓe�`�D4Rc��B*$���^.1�_:u�@ZQ�4�@$����C�i�\2�J��Z��+�Mf��L�ļ%��d�a�f�z'[��G�M;��Mh�n��=| �2J1�l�s��jg[ Z��+z��ױ?B�V(� Xj�扂�x�jGeIt�
�'Ñ�E���+]4�J���`��
�,��Y�B�t��K�������,��9u�0{p�U����%2�GL��5⑹+U��ջ1H�N5ힲ'|x�W����AXlxVHYEB     896     280�V��.1��oъ��*��x�|��!(W��`��4!�|�b.�A`��::�9eyvdt
���]Ra.XQ�N�w��p��²�Յ<-�s&E�����b�\��.^}��V�s�|ً�R�=����.X(��v��KMSt����Y��D� �Lf�y�͒������P�Y�r�?����]�f_X����1U+�%ܨ�L:�sU/O�j#���A8��9�dUl@�N0�9�'��X?��diU]4;��7��y.%��]��F�wν��]���d���3�rC���V��zv�Y�"<��>�o_�lW���'qu��&~0�*`kh�%�^6�l�#Q�L��6��O�  ^����Y���O��E�\;��w���G�W�or�����k�AO'��i^�K��2��/�]!������fH7�n ��4 ,@�"�T|��A�v�%Z�L
�@;�2� ���C�Lsǒ�F>+�����־1m���:�·�h�A��7�M!�ك���<L�`�I*���<Š��,�2������ $F_k��Y�e�bf��0vi����X�I��y�����e��p�$�)W:tﱀΐc����}��Gڬ�?L��P!���2�A�