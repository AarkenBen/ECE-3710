XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��vQ^Ʋz��\L;P���ߜ�� I��	�h3G�e帕 -�[��Ȉ�8=d�~��/h<�84��S(H��� �(u�EʥN��l�2 �j.��?ru)�.���"������hZ�kq��g���IG�?��Uc`��^CБ��+z�h8ZqהX��ʀ^@�E�g=���]c�
�T�ݾ��,�Y���%&�wCG��Uc���,C�h�G)z�o��$2(t�dAq{[��a���I|V�j�������������`]/�}S�!����h[Zxg��0�<�J6�Sk�@�=�d�>_�ro�Ee�B1�n&Iy4���C2�/5��'�k�a_;N��1�T�A�����H*/����jJ�M&ݞ�Kau�'�*��4o���"]������:�!TC��(	W#�p:Ą��L�e�rqV���l~Qu�u~��V�\�\�և�a�`2��P����ݾ��ʟ5C4�˽/�o0C��n�)��b�����P��!E�,�B"D�Aq�
��dn��PWc���������=�bΞ����G�=���=ĭ�^�U����I�$D�m��O��y1������$���Ճ��`I�X��|;y�t6���ݻ��jiP��N���C��2I"�( �tay��(߇��BGx,��_�1�
b}��e���	�Z�����mٓSd:�ԒB��J$�)����5��P��v�1��o=�}Sq�� :�Q�K\X��p����{! ��Y�=����%��t7XlxVHYEB    162c     850b���m��M�!w���l�~�����<��#V��v��i�O���E�G���?���#b?�˱��y(+���0���9Z+`�	}LSJ>�5|�)�����q�?j!�/J<�`�9�[ye��� %U��x�0����v�@d\���-qX�U�����"�Y��2o��c�:��P����N	8��t8Q�a�����nN�z�!��]C�hsD���uT:�E�v?�3!�$�C<�%�W�j�+�>p�%���ٵ=�E����-�Qm.3�d�A��@��g;�X&�ރf�,��HZ�Y 0m�*b �?����8&�UQ:L��V=_A��-��i�@i�F^f=�y�c�9p�8��\��A;�[��S;�]X�P�ص4.���P1�T�q}<�4���9��vD4l`��ፃL����4��d����_�x�<�e�f&\!�h?{ʑ����6����	3EO�i
�s�^|��L(��:9�6x%|��=,�������z�㊭� '�kߙf�r�O!� �m��t\�(M�W�,4�ft���l�zLϼ���
�X2uA��T��_�B\;�h�J6�f�;G�����~�PFQ��P���񕋑�=:F��G�q�w�G;��c��X?���z#9�t
[7��@��f�!�
�z���O�hAe�}��ԭ��"�Ł������a�"Ju�RL�9q~��-5����jg�SD�X=�f;ư��w5�w�����H%w�׼�Q=>�G�8n���u��㶤mγs���*�G}���U��%��k���˰��Nrd\%�g��X�����'?'�S�E �@kp��;,��<��[�p��R�~94=��;�d��"�N���(f�
�AS���/��\7	-E� ��p�&�O�PN�K{�n�s�������޾��N�����9��h�y��I�,H�?�L��(TN��L�H�� j��$cF���O5RĀ��\N[_�E?b�q�����7	���?��+FT ����;�6�p�3��h�~�m�V��;0<ۘ9a�j�T����i���֋����ǑV���h�дC8P�Ĥ����#���Md��E<{�ͼB�Ac����X�� aQbhR����z��������7�7/�����ɓ)�CAP-��qHA*�'�ip�$�Ğ��Rc�lc���[t��HQ���t��~�k�|0���d����c��(yZ�K��U�qp�+X�m
#V�2��+�Vر!��0>�e�ƕj@����z�:pVoXh�2<��Չa1�f�,�~��~�z<��Qo�؏'��9A��(��7Z�8����=�=O��	�ڸ�"6����y�35�L��2��8m���U?z�hj��o���H�vLc+��|ᬦwE�T!�m'˶��P֐�����v�6T_Ic���7�Y�>�c�;���q�g�r�+ߍāy,7�d8`�&~�H·�8{�/K���!@�lz��[�縂�Ǧqy�\݊5r�r�uz)�P5�S2�?��9Q&iE �1ڐ��5l(���5��1>�|y�)*'����.	�l�A��^8��j�T1�.���Ojy��&�� �GNڋ�[�3���\X7� �y��������4�흺����A\n͂��"�K���H�����IO��}W���6��*�3�+��*�X9����^�ӷ]�c����l�D�Ru����f%�h8�E�syǽ׸�I)u�k=,TH��H��}[8�m˶�Ϗ�@4�6�
���"��~6bMO�^p�)Ͷ�&�\��2�|q*#���[�i�ľ~�0�o�厖����WA���[A��Lg"�:�]�4,�1+��5����
�? �t�£t�2�h5��mD���3��;��x�ׂF�
i��!���BQ�B�a��!���߻:�XK�S��_�׼D���.����^�����l3�	Ϋ�ɪ[�C�z��N�߿���s�t�ڋ�$�td���c�����1:�������p��
g���P�L	u��u7�u*������}gu�rx�f$B��H���|�$҃^:��'^�H��5�p