XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n�Ҡp���{�n��*��t�7�]M_A�ՓkB���",��$�AҰZL���i��U�3��F��y��	��(a�7� *`3���� ����Be3�+�B�n3ǝ����i�5���ǚ��-�%�ހ�B��{���K}l���;&����s�94X��,���&b������ �ʻ�e����F&Ɂ�����O
�����Bh���R�������ҳ�t�H���K����i���^��U�H�����weo"q�������:A{��L2O�O�/h�P�ݬv���8b��4V}"G{�]�nD�,>w�+b'JU~����!�T7�ܢ����7�keZ	=��V+:�������������B�B�Z��Ay8�O tW�
	��pRf��l���ok�?���q52�\��Y��\�|�?\�$'�L1r;��%/S��6�����Jx� Ӏ�e����ͤ���X��>m��>��?�(8�\Oy�J�xsu��V�`�-�7M�zh����1��LW�i�r�"E~��u���F������Nq4�q��?���m�(����<��Ra����>&���K�S���\���J�rA�Q^hח/�<����	Q ���m(KM���ws�v���e��)vV�~Gr��S���Eތ{R��g����m?"�=��wMW ���x#JeA��R�ͥ"^�*����w ��dO��`$���;��
ڭ�iپ��so��D�%ѢXlxVHYEB    fa00    2950AOV�[�&��fKF��8>�'��(c�ĉ�&�Iw��ih���!µ�qNT��R[�B񦯘�1��'jKG+q���򡿘��n��l�e����T�J-F�j�^=\�9H��G[��J[U��է���]<�I]�sg��>?�و�>(-�~'E�Le��ʭQE��w.�2T ���Ρ���Y�������8�d�<�-�3kz���?L�*98>����.�Ѣj�Ǉ��b4�^�惍iE����g��#���8�
N��щ���B�����0�,��Q���4�K
F��J7\�娐U���Z�ʜ� �d�Wfd��n�L�^Xrڧν~��c})��
��_�+�H�4�7�
���
h�y__�5&���0#%�!Y�'���p~혹��WV�+Ba�w�*3ְ�m܎��-jh�?8���48���\sG�����5�`���7x�x�Y�3�.!!�YD"&��s�1���xo�.Af�۱�/��㨲��)�ō#���T���g3q��Aa����@�xN�a3)�H��P	&�r��ƙF�+��8D���cO�����ܷ�|+8�
�3w�t�>f����bݨ��F���ˆf�6������ꇙ�<1<�ٜ;�w�T�?�!�&����$���/�}Lp
z��M�[���L�� 8tR�u V����[Rb"F�
D��Cj[��.�`5}��R�ҫ.�Jn���e��BF��l�=�#�a�4Q���sB�h�=����F��;i���}*�����`��'k� �yX5�@}����'d��?OǅҋdS&����ɔV�}~�_���8@0�c�"z�lH��_$�(�X�� �1#`g*��&'��{T!k�d�w�I�̈́-G!O�jc���8�
�L���O6��p��X�xGf �
t+S����4G���Z�-�诠I��������މ�$4;���p��9�ς��EN������>�/��q��h�]�8��cLL$C��b��Q@�>@�=X%�G)�W�ڑl�z9�[���<x�v���zjO�m_BW�	g"{$B��*`�ok��L]��`^�UHʩ����V��)��ٰ��i�$���6(K�}��ðA�"��p��*�}�m�W7^�E���y{ۏ��EĄ@cT\��B���? "$	��`�c�'�1<���GoA��~�%1��]ȯ�	T}�2]����S@PeJsW�����q��C�f�>���r�G��p�5g��l��OLi�W7�ƞ����&O�xO��K_E�(�'�o]�#�?f&n�j�է��Y���I����~�!k'X'ß�f�2�QZ���C��S��t��6�7���ܐ����FF��w�����
}�{<'��Ah�N*n��~4�x�[��Ovτ(W��qN����K�+�0-�&݂)�����n)���BY����P	�+��ӵ�O���F�N���X�|�M�!�::��p���T��:����q��ٽ����h�X�s���gd�za-��I^Cf�����*I���D��$#�%��L<^f䚦Tl7⇀#�[W1W��w�C�!�C�}s��n�b��:��cCƻg=kų��h������dq��tW
�wK���j�"����ư��G�۵G�9�PZ��p���zV11&�H�x�F�v1<
̦UՔ�)"�4VSc�~0:zN�M;!��'�S���o���-L�G�ō�&�,�/4PHtz��⇖�g��"ǝ�{w�M��T�?��+��>r�~���FVJ���ύM�����䥽�w�n#�1f5��n�'B�5�Q (f$.Ѫ&j6����Z���s,a#M��f���mu�C�+�I�pX�z2���{��!�-�����Lw�-d��d���) J�dǲ����}a����즉�,4�p���#;��G�UY��[�5����8S�K���~C���
��8J�J{��МE�������53�Iżn�!���C,g��:	�Q~�a��k1	?_���~�лc�ͺ�K���hs���A���t���tU����ϔVL�A0Fm�,%��#���5`�=�Q�_�hbqI&o�Ǵ@��3"&�����愱������aVOt
�Z��}2�n,��'�	S�*�e�}c�����y�%UzA�M��Z�?�h�e���K�bE�"��N��ɏGe|Ka����3vP�l�������'�Ѹ�L��P�$��h0ٮ����-���׭�ۯ���_�ð#]UC��侢X��+�熧>�Y���W�8�)|�̂�j�2���;v�B���:Lg�vl��^�p0ڋ�D):-��f�3��e�]��dASWf���N��f�H�#ZQ95�4����E5cK��.���5��S���&n�_���mɃ����D>v�b�$��a�"i�5�w��QtV�f�t�t��J�'���`��O#����Ҩw���� ����t��R�6����`_[���o3�̪Dx��`��`i�T��A=�8z��+w�H��.^�L	9򉦁 �:�qp.���8���θ�G\�]A����k{�v.�숀ٟ��V��sֱ ��5����p���F�@���i�]IN!�vJ�aP�9Ϗ�!�̡;g��3~��zHH[��R賤�!��)�T��U r�#� ]u^�,HH�=tڬ^B�t����V�!bo	��	���F�,�H!�Y$I��	Hw&��,LFp���+3�a��wbb����Z��ҹ�z�{�D"�=��Z�����S�ː(�Yf,T�����i��x[���k&Ў��k>&%���|b|�Г��p�1���ylן�[;�d3���fR~x��j������ ��p�%����5��#����I�VE�q�R�9I-���|�3W�V�"9�lp��um�-Y������i�9�` Z��0�C�j��M(����j:i�(�8�_�人�t���s��7�S�$����u	Y?���2<��3�%j�V��]��g/�V�!}����ec"�%-f1� ,%%�돠^`��ȵ�H���O����pfHٞ����)$����ǝ�'���5f�K���&!�[7�U,1��B�����Fc�E��{.�~���%K�y�"�%�t,�ļs�v���˷b���\��9JYW*�k��K��c��[�b2��P��e�pƽ�� ��d�o���� ���!,+��`	��9)I���KɃ�p�ڰ���(�>��L�R{Ӵd�r�C��6h��C'=N���l�x����d��n��[���TJ�;X���g�p�:
i�=�����E%�qAp]i���7�U�'�{�ҡ�*G�t�7�{��u�-��Z��w.����a�:V-y���փ3_!�A��6�n�	�Ɓ��S�_���Y
`�O[^P����Z���W��c5?ʡ*z�;��5#Ns)���T0b?��ru���z��>V�8�����ZT��}h�d�D��h�s�����!Է�����#3AQ��?�b��#�#U�p������'}��J��	�s�ު�-fÓv%��(�mU����jV��0�s��}d����c���F����U����w�C��Q�n6"餅!v*ajjW+	�!Ր|Rz�}�\��ȮW9�0���6�TTYbA}2H�O�>�	u�
�r��!�@{4��t��,Ha5	V���R��\x��֑���9|��	�΀^nm���A�S�rs���VO���ꏭ�ڏ[f����W�||s�Ǽ��V��aB�C�@���x:}�	�W�$��3�Y�3�� x6�D;�g�P�;�3��OK�~���V��x���>�d��x��;�E���eo���8ذY�z=����ƕ��V2��>)�����Y|���0��_hrdC^���B'�u%bU�IL����
�[�C,O��
��p���R��I?�O��	|��+�52(������+�����:����n�&��|�EQ�_��Jy�̐�d���ډ3��eW��8G���������+k��\y���j�ޕ�	+��O��X��9?�m!��}ڝK���闯i�s�n&t��pc�������iԨ��ŕ�
��0J֌,�����ϵl`PNn�v�?^5D����g�ح*�������3���zϦ�}���� ���=���f����L�/%bd��,�/_�Uu(ƻxl�cxz���Q��t�@ߍR��_�Ʉq+�(�@�����j�?���HUԂ;�b��Y��e��� ����*~���\��������K!3~2����v�^)�W-�y/6���V�/</��j�+!�$4`��C��y��3%�|�zQb�\8g)�K} N���Q�ϋ�ɯ���A��c��_>��x�ݱ������c��������~� P�[��oN�y"mH����B��d�^��M�:�{-�?��������1�~`d�P�������<o��N|����*'���;��N/fX�����;��N��Q��H���ϔM*�c�!�i{��n�
`z0c�g�Q��t^�kM�1��W��@���7;=�����~H�ōq�X�_�Q�}��ǌ����Ni�ow�ü�����X�(Bu�y^��^'g@���h=P:��Y��8Nj�=Ö&�=�:J�t|4�3м��_����� �G7K����AP�-�jSb`*�r:;����R����̠�_�3�E�k�P*�~$����~D��W�a7��#;7?��/�?�K�Q~�h��rQ$Z���wS�^�C��`YA&'�9��Ȇ>fz�c-� މ�j'&媏�����R����Aל�� ���G�sf�Oȵ6�,�1��y���5S��f	p�_��g\��E��
]何Re������ {b�z�]i҇���X-���pT�e �� C�d�!`�@����E���J��x>qOT�ܹ@=�J�R�4�[�2���e�\>�۞�b/:[h66����G�����Y����W���v%��P*������i�����>��Anޛу�9������ՅZ}������������Aq�B�[�ڜ�TJ��|��I.��P����.��"bj"�z��e�`&l �,�[6�p2 �U&i]�Y��dM���
�L�������i�i�����h��aL)�'K,��Mm��m���̭���J�Ȍ��@\*�+5R��dkSt+/'k�?J`�Zp(� R�@�?����0���H����0���3�({�!���i�@H�vp�����K��#��M��(k���K7b	��K�z�.����:�٫"�� p�O�W�@���߭�c>^wy�M���V6\wZ��X����caE�)��_L��U
��ţN��x�)ҽX��|�i�5�GꞀ�W�'՟Da��?CХ����7�N��|m�˔�AL-�Λ�8՘�����`�|��$[�!i� ��]�NH&�c�VRQkmte4���K[=��d`�^3��O*3�P<t]x�Bǜ�*G��$�Q.!����K�:.:,�'ݔ|q����Ц ��Ӷl��y1O!�*��f�RbGB�A���}ׅ?}���	ԇ �������v*��r�gO:��E���a.˛��e�&���H$���Bv��Y�sI"m�*�L�nJ���4�o �bh\���*������2�Q�.QXC�P���~E�,%$�i�oK�4�K�7�!���uB���Av����C� 2��L�V�%I��Í�$��}���ڴ��q��4�cj�*	qP��R��|�i�4iݣi�V��7+{��	���V�*C�G(/r��8ޣ���?v����b�!���m��J	�@u#neE�M�Jݵ,@G��$��������d��E���(���2���t?,��X�W+���o5OVE��ؒ.�L`	'���Q��]����l�<��<=�ٿ��������C���jhc�����<H����I�'��σ��,X-�>���ɚL��Aj�~�%	�<Q�����͖�o ﵼ����~�%O>x=-�ru#�F��Z����+��;�w�`�i|�1�缕�B�6ٔ;�����&���o���nW�*� )�**o��v��s1H�"^�k�Cel}�~�E�� x�n���9��l�K�<��y����Mu������3(H��U�p1������wʼì&���
!�S7�h�~9��`��NP/���2�S��������7���el��a��S	,�A�l�hY@��`�� P'N�έv��F[�uj��sEY^�Ns��[&)�҅�μ!Q��Y���ǿ��ۈ�tsn� ��l��']�t^W��#����K���џ�5���U&#�q4�`k�]B�u��x�% ͦ�c�T��������osh��ɴ�<WaU]���K��*f��ڹ����͏��w�a]��6������S4�؄u���'�b��
�����oč�����l���h� ǧ�^#�{�3rq�uqX�B��mlDu�V������֐��M���yာF�j���Ew�K�>	)ߋv��v ��;(*��vݸʃ�	p�M����G�����\�G��auq����hH���`�zzeV��h�O?�ȟ�H3Z؎Xt.���)�!-\��Y�Z�{�' i���Jl���D?!���� ���j(�	�6t%KD�O���y�
s�aKDit)Y[�g�4 p�	�ó�0�%���]X�
���kɆ`Q�kl��wL [�;�gm#֥�;��ca#^Q�����8E�-y?
zb�c�c���.����a���Q��86$V1�4�t��M @4~�;��E��Z����Ю��W/f4[�i{� �#JK+i�OJ�z�n��-�:��(Ca�aTS�q���h� ��T��I\Q��v�8����?g0��_�!6��~�x�����|�K�t����C��q�sS���o��j�_NL`26���#��.�+��	g�
R.����1ڱ&#��أ�Т�����(�Y �*mb̠Ed]���(0�s����� J�ku�2����-����)$+4��3�=����ਫ��?��^���;�J��A_y�1�4��<3J&�k�m�qJ�_[�c�?�:^��-_��6s��*�uG�=�@������T ���O����b(�&I� S�|��au�/3G���3��硙���@OPD�f24Y�B1J�ã/��L�����E�$7��>�Vs��30��>B��(�I��Җ�&����*7��i^��ߨG�j iŋY��}�Nƺ�*���%�N_$�Ly����p5S���~�����L��#��Jn�V8��}�g�wu����G� ʵ��#���Շ]�c��4��n� i���j�	��V2�u߳Rp�H�}�� z�9��S=�r���G��8T�<B��щ?�"���cO��.G e��<�@*�ި��wD'��JȖL�������)�͙gKQ꿤��Y����(̰�z�VM;g�=+4 ?��8M�m��x����]����Qd}�9�A���sA'bP�k;smG-"Ø�Dżcݽ*`C���Rw[L\�MM.��$wW�4�p(~dyvG�v���m��>�H����)���Z�m8�v�*8�5�s��A����'E��k�ן���?�VR��t���]�zh�o�R�6	ϔ��椠�	<�W��w�-:4����뉗����7V�$�x�Yw�����C���j7{������S��14��N�17_�=e;Cw���~���z�z��d�=�ڨ�>��55)$)P>ф��x)�sT6��U��6�p�j��D��:�C�� s�F``d�ɫ�(q�˔|�䷱^���3�N�h�)��Lꪥ������V;_��OG�ׅ�|�Ț )+��*p��f�3�%�ƫۍ|�ıc/(,����9,�*�X�I?$�r��1LS��+��H�E\�ԈUy���k T�t���U<)�|�ؠ��▯<���v��c
�y�����t�ɠ�{"��u)���x��^f������!,���T0�Ǧ��nJh����U��h�aq�]�i0�/,��&6��}�>�y�_H���O�\jc�� J����m��P��f&�N�ňH��B�(��B�P7+n�����u~O��v)v�{�,����X��ۖ�Ib��^�{��i����n���VY3�eD�76kȕ
H:���T,�ID�{&&�qO�ޑ�1)f)/����p{�lX�#D2;���\ְ�EW�n[�%r�Ͻ_~h} U�@���Ӈ�ŀZ�����g����~�}d抢������d]ɪ��|�'�:H���)DT�2�'��l"C�(�~�� v�e���!ǫh䮪Fe���'�c�6f"�ȋ�^��0>?�#g��4Ceq�!+|-E��������m�+�%ӿ��D<�8��"��=������YP��F��u��-� ���Z�]�Z�#�(oQ,�L�'��&tЂ�D{��]�ǣ����ٸ׿�;���R�Ļ�����wl���u�l����U:<q��r8~���10��5�����������g�"�2{�{�c���#j`�J怳Ew�v�˨.�1��j��p$}���UsN��`�-r���'�F���&
�q�x��upk3!̝<$!2��lDݮ�>�4��߅�Bh=珚#�Tä~k�6���]�Gw�g��lg'X����P�2Ұ���6ט��Q����Y�:3�\�\j��Ie!]��>je�6!�=�Ĥ��,C�L��u��Z�n���0��O����^����rA��aI�^s�T����m�_�Ñ}�>oJTY,b����MV�d�e�? H���2G�?��4D+B^%��n���� ������:�+1�:/4J��O2m�(�o�l_Pt��m�4���N%M�"]����a� '��!=��`�m�O[~cOo]�s�Ώ��uγ���P�CѠr�U~)�� ��z�I���[�.r��.�*�^+g��C �`�-a��S�kj�w6��⯷~z��R�n0CN���0n��E5�¿aN��_���&��lZB�i�`�'�����'�M3������3�3����*�� �ҌPTȶ���c�� �M5.O��CQ���v�I�\��T�t�Qe�ȁ��N[�MR'��U�L��$X�U�WI���s�Z��]�,�i]�(;�>�z��� M���ya��aB��7��SIT�s˘��X�}���x���v1j�|3f�\U��p{-��ٖ���j�ۓ_���W���?r��<P�M�-ڲDą�oL$]���dR�V3�����J��[��s�I��ѧs��쫈��Q�[�y�{�9���_l̝�8(6ɾ�P;�/�E|3g�e6��N�]���"ˎ�\�3�8��Op��q���욠mе�]m��K���L~�o��&k�NF��j�?�ζ�K�#
�y�e�pl�l�x:>�OУ>m2d� ��SBpO���O�����0�4L�P�ȴo�����7���ղ��_L3�s�O��j��5�"����'�
�$�1�_U��"䷂�8������q{h9R?y͝bN�$�x\��V8��$q��&�B�h��QR��TܹH�����;J��=� [�����H�+�d�z���o�e*s��KckK�����i�aFZtM�6Opr��.Ƿ��I�j��=U���^;��s�y�w�_}�[��*16�Aj�뗓�m��%�vջ�s]^��a}��=D�mP�?��oV�օ�1
J�H�Z6`>mOB��J�>��u'���խS�,B4i�	o��gh����o�9��b6��R�Ɲ�~�c����AAc���)���EnUV���ڜhk��������$N����3��e=�c�R��y�<Ʃ���"oʇ)B��D6q=XY��2���B�=`��3	�-����@�6!��S�?wOsF��j2�mj$�{�U�׶��ůc�������:�����j���wg0s�`�=$0��l���
��n&����K뀄���Pyŕj#�}�:��@(��ɱ$��x��v��F��=���_�W:e�	�Dq��+=���mD�x;$j�� :��WFA$�_}4���U\�-�������K9Ʃp^�����iF/L�\�{8qu =9^"X+�y85���Ru"1�K�7r��־���k�q(�ǎc�)��r�*پ��1PP��CS]𶃐���c��p��a�Z��hI7��g_��V��5h*��>�E>������&�̞�U����#��'��XlxVHYEB    fa00    1e30� �2���$˸۱������Jy_z�%���éf�i�Y�jq�@�֭���VMzf��W�Jw�x�]$��D�|0���3h�=%j}��m�!C��f�5^�-��`"�$��_�ۥ�nw��& ��%ۮF�H`�-���p;'��w&������X�p��P�Do���:ظ��D���~E�BM
x���l���;�ۡk
0�EJ���H��i��;���R�dM�Z9S�o��a�hd�D��"�£�`�?�Rg�͹ix����B���| >��8G�n�1����c%�۸H�����֑��)�D�84��iz�;�b���޻4�ToY�Z��joM��	xY�ʸTd�fܟZ�Irp\�!%�Wx�ȼ�d���i�:�K:��BP���������0$w{y'���Ŀ����cGy�S���hNC�<��F��j��L$�w;R�߷9�.���4�����H�'7���l2��O'�>-���%KE�ѣ�A�zRPGK�2�3O�P3��v!��(H�t����t���yY��N��S����9�c�D=����7����� �Du
�GO2-��$f�5�̫�>�!�<�#��f����K�H��1!HX�UC(��Zh�K���L3�mg�(����xL8x����,��4�e�~���Y�ݼ���蒕�����Vݐ��l�¢<��9�8��Oi����­�?����x��q\t!H*��|�%h7��]�5]d��:֦݁���:��(s��hJL���׶Qm�MRf��Te;\+"/�E��-䒇���<S��}bD8���;�(-р5n<�1��h���/��4_`P;}Ufp�L�{�@��6�p���L�	y���W��Td���]n � ���B�8����� 1
�3e�~�ݮ��&�����q徬�ہ�N�V�?�ɿV�[������˝�%�6j��H3��k�`��p�}BHX%ُ�N�����Mv0s��E�2��R�`]hf9��`�[�j����tUK�?�I�i�j�D� ?@���lQU�,0�h�p��G��� �K�/�/=;�r'h����J�3��XMʫ���#�]l��c�����*�p.�0���@�Z��r����������V_���Y �{��(ޟ�`	+�'���	]_���|���_��p)�ģ�1z
��w�T�����D0��Д!͵ 苉Ĉ,�Db�S.��Z�<��#.�4�@���g��
R	̲M��SEN+�f�F��P��( ���wOYW�3�
~�"r��A����l�C��R��`���Uǡ:���;Pt����3��`R!��M���śU����Yf2�U]��x�E7�z#1e�;ͽ�xHT,#5���磹֕��y"�I4D4>�-��6]��$IUwY̸a��V@�U5�)f��u�5Ɓ�oצ~��zȈ.7�q2Ґيz��i��W�+���o``����e�g�o7|Qa~:�;�<�W*�c�ǲ7b�������rB�����]�P��u���b����l H�C�丧I�䵌�i g`��%�O�j�.��)�-�&�֫�}:;ju���ōD�ꦈ_n�j�nL>:>���KL�z#{B���a�d64˦�{�|��8dU@x��n&Wf.t��(��"Θ���'s�O׽����l��ۼ�ʎ���@�վ�&�d���}��7F h�A`�cf�0��{��LY7&ro�5h�%s��ډ�r�����K�)���R{�@����\���Kƽt8���
���=m cQCi D�ya��A�Fcl�Ie�CX!�W.��[N"B.!{�1��h�C�;Cd���sj`�'��%U�����V�ƍ�©�!���p\�ٷ<��̜��[�L��7%M���9�����G������E��@�oj�&� �d��ƢlN���ꔓ� /.�&,~�Y��c��o� 	��xR�<>D��6K�K'V������}O��V8�Q.�_�i{˄���:W��p凨Q��a�d�	Nͻȹ�fN\��Օ��}�O��T��b{�����|G���ķ��	�ʣ�b�@o�Xa+?1>���:�����7�T�'�B���1���������1���)�uf����A'��NU����!��J��,�,�gc�*�
Q�U�����l����p������J�+�Z��P�@����6��#,�dB�KSख�k�$���^�:0hP+�>՝�sp����q������������@+s�`&�l#��a��� �-8U�kP�BB�
�<Ll�������4�x�}NL��Q(#�����\�*���]�SDyC_���(��y�����[5��x���W&��D�d9��
�Ű�[�?a݁�ո7��wjulf`�+����׺
%)�ض�=���ꂂNY���8�@F��."�}.F}$��EV����Q�ys�l
T��6�P٭���F.�u�AI�Ơ�S#��?����8)j��-�1cSF�?�R�:�+��[6�9H�/���e;޷�A��(����l\g�dnl���y�"��:�"�`eV쾗Q�k��c�a饫{�K~�N�uK,���I��}��Oqn%}iQby��P�p���H�et�1������{r _�!M����&��ޛ���q���]�L�-{b�׀���1 �q�/[��'*49m�����ȡ�%�5/�_Y�������XE�ɤ�n�NY�t�!��V	���KE�-���=�i_F,��Z Td�	W����)�y*������|�6��_o����¡�w¶�d>O��?b�Ie�r�Q|�Q70L�E���wqٚ4o�2���3{��3��力@f�/���؉����&�2�I��A�,������>�K�WW�;�������@���2L��8�j�l�P|�p����v�J�[	�R;0b��\�>������%�B��.�na�u0&'3�J+���e���G?ptY$U5[Y�����W ��a�^*/��E0[���w�a�LS�}��edh�'�0�
�}�0~�V���[m��'��]�I���ڴ�;��.cտ}�f �W��숮��?�ŀ�?O���=#3��Tf:�L��8�������I�%�)����~ӵ-�"U�Q�B]>��aAt���L�]�b&�����@��]�'Nߠ��V�r2��o�k�3��'��`M��?�%�:�j��G�㌌�x��Y��b��b����.G:3RK��� VU$�41a�ſb����N0{?^�]�[(Z@qu��"���b����/��wD���X����~��-�T�8�m�8����Zd�9�G���H��p�[���i�W`�,`�����ywiX}HB�\�-3�ِ!�����ɼ��B�l�/�����Ym��^j�ժ��N҃�<���������?_3�%Z[��^N"�{'�L*��F͛_-�R�݌ ��<Zo����Q�..اg.)���?7o�����Dw'ۈX���Gtk��Vt�
o2r+3�5�E�����'�?�����"����>������]�7�}��)˴��`��}�Y���J2[ ����i�v��N0x��S>O`Z �=<i�Z!��ӆ�o���Qv�)O��I��L}�;o��=����]�{�`E��9�C.�h�_K;晨`��tj��J�1���q'��/�D��t���ϣ��9�� Cf5��摄���������g�i�	�j[z�ĪN�Yz[4g��`�o����p��T��MX�w��r�&ˎ�1��<�ɤ��B \k^�;��5\Yg]ɟ_����O_Il�E��Š���΀ �yW��Ff,x�j�ʽ1���38���7��KOS�Μ�j�'����e�o�|�K)f��V�p�*��HZ񓍯��A�Ã�@֨��̃�k�u:>�g�rk����|u,���C�2���n�tȮ�`�*���9@p@�M�����瞧wGO$VE�X)��H��J 6�1*9������<>i�����N��49�	n}M��h�\ڨ�9jrƱ���D҈X⢸��Q�}L�-<R.�h�l�w`l�S� �ȑ)��5#$�r�����y�x�T�Hn�$����f˘�����_ˀ	q�PK��}�~lOEB���ay�����V�	�+K���:�y�"Kc��u�����$#��b]Dj+澴Vnf�ׇ�t�]�:�r�iƒr�Ζ)���wu��ƚޅ	�u0� ~��R��?���F��iM��X��i�(����j�0��"��N����~&�֌��a*��ᶾ��Go���U�f"Kŏ�&�ܖ��YS�Qn4����i���2ht�&q;�˳&Ƭ�y �Ý�	��I����sz|����9��̚$P킂�Hl��O��Z�*�� G�{�#v��ݖXd'�vx��{5^�+�9��ڍ�0�!}�x��'(ˎJ��t,�ii܅�~�%� Jn��֑۽��+Jf�GU����`�f��]P�S�r>�C]�ա�UL;o�<�\3��`sv�����_�J�
�&s>�ᵽmR8���Iz����D���z$���Q���9��)���ԗmK�?{��%7�����2���xգHh��Ngcis��PI�����3����FQ?�Ί�2�olAB�:� ���/+�2���!�?>r[{�����q{�^3-���c�Ȟ�l6���ٙ�W"�y��Qd殣g����?1@'���+ؖ��W���[��:^q��D����e�1'Sm���Q^���u5a<�a�x˂�l~-7�\�ڷ��^i,n_�o��j,��}ʋf������;�zL\���]ug����I������_�A]�> �y�Q�äۓ�Ԥ&j{K�L++6����T��ݷ�����f)A׷��`����v�����LAY�^7��@h2[��#��l��K��!��բ��p��v[>�p��_ɸ:?AW��C�c� �t���*],�-�Nu��N��|f��~r-���w.$�A%r��M)�����x��1����8�����Ϫ�Q�!.{�˿tG�IԄk�ƭ�ămE�qU/��6r��p��ό���?�%�lҞ���`koh�����2�@�9���Slzg��^\0�tސ}Xվ}�sU!ea�����"G�ܼ�=��%�"�/��A��i��5�'�"bLF(�;��4_atU�Ԍ���h���O:�NڞԜʘh�7�L&�[Yܵ�w�zR�O5��)G��;\bw��w�2LA�n�Kԉ�~�v��{��SAݘp�k*�J���p�l/���Z�ĺW����嵈�
VЧ���@h0���,s�H���SCnBoQ�b�����˧��,�E�A"C��\,>�?�C��=�O艬�d?^�W[A��8�rm�F��u��T����
�XN�����M��nfVD���8gK�l<�۽诔e�����a�&�V��#�,ֲ��.�4��ʕ��y���J;�EС��3?4q�
��9r����y$�!.*p��	�0�U��x`�������UJ�#���qAr���S�b����6�
/u'8��w��6܍�[�J�u ��7�8��
����m�F�74|#�W5#�0pF��ռ��ǷzX��s'�?j����y��o���VXƪ���d�*MQՎ"����^`/�� t� �̑�e���@0;�Ƀ��1~Eʿ�2z��t�urh,&�F:��V���h�� :�r����bս�nE�q%����V�o��T)�F�n*Zt��;ֵ�!Cx��.��I״��`hZ�u���[��;;F�o�܌X���n���^��|�A��vRL��b�d��%DLk���ҘƂ�@�;�6�h����ݎ��D�P7��a�����U��Þ7zkxlf�\٥��ԏ蛠t�Y[-�h���?I�f�i��Ͷ���l�9�8Dh/��c��qeT���#�?��'~��]�߈���B��5v;n�׊���g�s4�s�lZ�u}G���=S6֫0�gxP�-���F� ��JP[������]�"��k���"��X-߸�=-��#LLW��Gs`	�NAD�	�1���z��A)&^AU���<�6�p���u�OZ��� ���؂k&XIJ-՗	�@H��&��h�$�OA����L�x��=�%P�.Q�H�q������e�B�\�ԹS��.�/���[����ב^/���*N�a��*������TzA�n[ QtQr������t.�o����w����	��L�rЕ
?�W��	�c}#�N�/��E���On����=S�ׇԺXyJ|J��=oK�^����6���d4Q�e����Վ�)8¢�Y��.�bVۃ�	�ɕ#8��W�1L� �ZB/����Sٮm4�����`[�
n��R�1�?�����&���	S86�9��@�%?�N��#�$ЪRNIҫe~���t���*�c��y��+^�%گUT�Co�`�׸��s�Ğ���޷k�eM���T����
�S�b�t� FF�YG@	I8�{����)~2d���$�nz��l�|�Y����s�E(�n\u(8����0�)d>>i\��zy���fn� ��)*U-���Z�+�fp�ǧ���g�L{���]ȅAR<qRJ�AAPU�W?O�3!A�����&\^��ң1�Y�sk�Uh��5�{�,��y�9��|ȡ�~L@�k�1.(�sNS7�7��u�l���\�,Ý�-���7����㊡��ִv�]��)2-Q0�.݆6��;-+s��W
�"#��'����6��4��s�6�Ha�3����~�����ٔ����Eɝ�b���.߆���AtS(�1)���0;�x� gאj��5�k�kK�f������F(?�r�#8������	C�`��N(=&��VMҰQ�x�2 �1�5b>$s��Z�ܞ2�p
�r�Tb���|nj}�jYЂ٠d'[|+�ZM¢��(}�^�va��<��%�L�3��M�$yCz�׭��̎��@/��|~-����9ߚ��s�i�[��V��vtk��^�0���st�L�jW/LPVw�-<�y\[W ]G 1���E�������{]� zv9�U	m>Q�3���肽ڸ��&"����XD� NԨ��]�B��W��)ƥ#5����S5s'���e��8^	��d�FaO�L�Ό_���|,sg,�˟��V�N"L[|??�Y�'XR��/��I��h0���W�H���4Zc�%��ʩ���C���#UXfғ�Q,tBwZ�qG$���s�V���L16��AT3A�Ϧf������A��rb��v
O�v��!�֬$�y���%�;<��R� ��@$j"K���m�w�z"`$��|�B��h����� y�7Q`~"����0z��>V$�Y�u�����F>M�n��_+�D���U#n�n�#2��C�a�u�̡�.�����&秩���!��؋�H�WQ�nӒWSR�M%��%����s�]H �.=��_���f�"�2EC�j'\����	|d�&�XlxVHYEB    fa00    1d20^땮�ڱ{�ԅ����a��Sgz6�����#_~�ٿЃՑA��e���nѕ�֩��<����F��@��MKb�,"�Q�R	᳋_�`�Z�J�ء�[}�3�ww�p�T����f��r���=Ր8�F�,�V>�͐6Qi�]��<�Z.���ٙ#��S��Xɷ��z��g&��)'��ը'4b�{9�zt�>*�$��6\'��E����bu��O��'b��z΋} ���%WK�i~��%I�~�U,�. 4@CC=�J<�&�� ��3�1� �(�'��ο>��uQ}O�m�����2|�S�,*�㸘:��;>4^X���A6)(�����15�LIQ*�e�����k��L��[P��@��D�$��Wk#�}���7;݌|��#w8=�u�TS�"a��2�һW�U��
Ә�(T�5�(#����6�:B�M��y	O9%�����S�9w��_ 0)��랱��4P�&�9t�ƦU��_���2�V��	����9��g�eѯ��lY�I{�Ȟ�M�#i�@��_��zq�}<�N���jAC��/���{��s������e�]��K�	��� �.��h�	KZG]_�Z8�&�1ip�ј�fXE��^���1��!���5�`��7���oH���+��H*$��t�ß���X�,�E��dH��zn��QtH��CX��3�S{*��"ss�$ {��^˜�Jҩ��ɁSȮp{����Y+�R�v*;���03�S#���7�
�'C�� ��R��Q�s��&z�/���|v�T�
k��w��kYl�s�s4��wy2"dU1s45�Oc[�u6���c��ɼ`�ת)��%>���1zfTd�����Z@:�	�M( �k�ܞ�����MO�!-o6�bKJ����b��pdR�Wf� �C�B�����:����N����k���'()q�t�唁Ϻ���{El&��Ǐ�h_��j(쥭��U�@/7b�]l��3���	:w�=l��i��`��U�mjt����/*~�P���_"�N��zQ��%u�s��I ����F�}m���T�I�)o�scHD��P�����b%'�6v�$ir�m�K�<ghU��a�B2��	�j�M�G���Y8��S�;�Y����)>2,]�	�$�o5�!D��pv^��P��?�׷�6sLV!f27wwb�+^��X�	��c)f�N��i���n�Z����،d￦/��	exRЎ��NY�1ahZ�O�A~�����j�[h������C���S�):-����Oa ��M�b�I?z�TN:��"�O ��/� ���e�/�����K�!5sD�A��}9<��Q��67����w|֘��+�@m�+^������V\Kj��]'��+�\��<�F��T�hU�՛����`�~��y�9�1��(5IS:�վ�t�@lO`A��aecpŘ�F��R9S�p���ǣE<�Y���ފ��=��3��褔s��,�
���2�=����5֟s*}��1��\�l���ߕ��z]����`���mv�����#�#y��_E��[賳�r��}�s9go�r6�
�s�/��vm�m.
�Z�+�����[g��Q_r�
0�s��>��u�g�Y�,��>Mnf�t4گjY���a�����yQ�e���_v��L�𲟜)#srb�죊Wp����n)�ּIӅ!��9�/3R*�X�'��
�+���0GQ�p�r
?�	B���-�R_ٙP\aj8��{�t���Ur@���Ól�o�����I4H���u;Dɒ� �F����GK���d��"�B��`�CĞ���s�9��Gj�8ݚ�JxyR��{�
�~P�|:�T+h%��S�r���3:���S��h(����=<��z�:2`jǮ@V�UG����ԭ��1��&.��d-��0�`�͇k�������4��O��2��_������#�@g�����|���l_�v���ЪO$����Fl֯�@'B����d��)���'a:LPoN,�i'����ұƢ�X,���!ߜ��$PL�}�C�)�	���>/��>�r;�&[��<�Y?��m
�%93�V�IO6�̴qL�i�3o�饍)�^����?#�n��G���]B��[����t1�w�၏�a�.%n'�=���9� �jIT���A�N$�hBqϨ��(�pV�`;��U�X��N+�����$�<��ۧ甸s�a�m7���I1��7I�/}���2f��������ԫ�B��e�4����ʀ��'_����R�5 �mڐQj��rV�Ȼ�A���*��9���v�1X�K�T�Bt�܂((��d!�sP���S�G�d������v(o��P[�?Xo�S8����eɆa�h�ۢm��յ"�ԋXN�U��x���N/C}N��U������K٧�hV"�@�QR6��f�I��ކ��,ұ�L�=���i]@�'9��Vi;�^6�~GZ�t+ƞ;�_��,�Q]',���.�{&/"�ܡlT�F�x�+�B�����g���T9M���y�z���'Xu�'搰�N
$��qť��8�'a�Х��{��r�i��Þ�����N>2�B`�E���a������o[�E}�( ��{ZF���~o�!#��&�u�v�?`d�h�����zSr�9��F�\v�q$N�)JWJT�Z�A&jr"�&�ÛVf��R!�{\���"�),�Й�5�H�j̵���{��x�hS;�#����h�t/�c�;Z_���W�,WR�������K^��d�y��󽲇�5�}��B�cI{@P=Y����Q��@w=d0|��!���8�M�M��-E��	lgt��&��j$�3k���b�����]|�G��Yjn�j`1w�Ѭp/���NN��إ�^�FM �3s>�xP���l�>������b+8��j�s�-�[ց7��؃����Pkm�+ C p�������5�	�V��Fe��ù�"�M{�mihē����»N�K��:LR3~�Oɼ�}��B�0�H(s�� zU-�v7 ��8A��X�Z�3v�{ؼ��L(Z���N�!����y������+�x�ceH�2�?��Z?;3Z u[mی���܀�[�:�t~�l�٨�S��� �#Ŏl��4	A[4�*xI�"�z�C����
�m�-�4��"E셚S��򜚭~��1)z�M�]�iI��P� �" ��0~��r���*�Y��,`W w�6����^�zr�]����	�f��/�P9,<�lʫ�Й���7c;�՘���VbTo1�=xX��ƪ�����5Wo��s�|�4˦��G���WZE]~S�g ���S��Ȳ+8��u��R�1��{/�E��k��tp(ƞT�ES� ��j,�ι��E~�p*f��
�9�
eB3����y����h#�R����}"d#�P(�M��_)����קպ;������i�8f˖.��9����\��v��_��#�_*�b@!���)d|�q�_�<,u�����ٍ�V#��=�y��	�a�����CJٜY�W�%E)�&Lxˬ�>\����ЯR>�p��@Wƞ�\I�\k��+�nM
tQ	�����W�NԄ(�(��^u�Tّk�?(C�1F�3_^L2��4��5J=��I��St�HTl9=q�Qt�\F�C��G�G�-K˚�KpTLi�*s��~���N�}��ۊ�]�������V8��X0���Qk.騩�G��lk���RbTf�׆C�����Ｖ�A�s/j~��!�����ڛC�#w���|��_|b��x\���l	�qm����1#����É|'��b,H�D��H��Ԙ���/B^NA��ͼ��}uU^�X���2�ű8:��^NА=k��W��;=�oL��]�M0v4�[�׀%��n�>G��ZvSS�v�ܣ��ǩ�����4�#
@��j�]�Ň��+�t8���ݣ_#�zj�񴡽�)����eׁ�R6��n�JX_��
�"l����ga0�'��9W��*fA�锒��n!K�ڽ�[=�-O����F3�~(���v��<,���CY)�J�0�=?��I�U%�U�Z8�Dy(�]D^f��d��	��FCr�;�S�f��~�r�Lm����☡�wF�"��^;5况�<�uo��T�TL��;~yv�'��k)?�a�f�kȟ�B��{Qx�~ �D��c��]i��G'�s��2p����Fj%a��On�wf���\A���Ŵ�/UuaM��Fȓ�q�7�Ԗ{4�+����,c<�.�|E�:O*)6�{2$��{eI�n>���϶8V��ˉӘ6!�R�׉�H�od��a�
c&N�G[$q;o��"=�.O�3�BE�&-��%W�8����@VnO�=�/s���zt`�bK���٨O���P������ �x0|xV z	�}�`w�Ɋ�0i�&�p5ο�L��E+Rh���7��s��$D��<-K����?���K�]�--�k���O��/J�TY��V"���r��ڋ��Q��$i��A0E�w��e<��[�d���C5��W�.��pRBA��p\t^^�	.`�9�H/�-���e�˧���m�,�!"cԀt����l�kO��0�BD/Rϕ
%�����d���1��~�T�4�ߵ��IGg��W���gE�z��|*�i������_�Nqx>�0��4Z坱F�V���$]Ih�*�ζ��وV/�D�����D�2��)���fքvcA(�s#����ID��2�j��Q�<�͗��V�_��+��VM�i�ҡO��F�c�vE��Y�l��(�� Yz�9�^�����%�����2�|*+g�ɝ��Z�uwZ�S�k�X~�����7�.�q�T=�Z���o��?Է�����mjxV�>�«�ȶ`�-
�$_��a����X{=�N	}��`\�[�8�˷��7���j�#H*�1��+���F����6$L%{A�%�Qt��2�Ex�gB��s����V@T���+�0&9{����L��#�����)x�F�u���h�d��穢���dtlS��f����sN�~�,��b�� V���|0d,8xOF���� L����+��R�t�:RQ_�b��I��a��'{U�XG��Iq�\o���Wk8+{$�.X�O� ��͓\�jM��]���;�	a��OA�h��zAo���<���x9�S!=d�n��?vNs!~7����z�eN��?K���{�A�Jo��h�C�7E������-��
m�/���O1��q�BP�|*���er��D^�>��p�Ӏ����]�S;YV�����G\��
גhҀ��vK�e�+b��Cy��s���"�Z���� I�J��Ff�w�eH��5�l�^�Ю
�i�Z�֠>kXX#(�E<� v�}5���c����0���[)��N��޵W�z;����Ƚ��w�"���f���3�J4�F.#��}{����>�	�rv�۶���R!�"%�0��O��z ˁSZ:�!���(؛7�)K0ݛR�p�58����r0�(�壀k=?c3�C�pI�	�� =����5���
sIm�u���n#����Ř0�L�DûI��y 7z����l��W�7�ht�	#~o�n���}�@^	vG��p�����M�1�~t���C�R�0�������9���3l;�[���@���7�k%C�m3�������7�b
:*H����z�Ͳ���I�l������`&;+y8����������p�|7�����MW�����FI9���_�-�m��4��]*��n�p�O�Q�Fy�]Yc��{;�h��$�G���B-ϊv�����z����D���T��)�6��K��u
Z\�5ޘ�_s�~��[�lA�z6�=����u� �zUp"?�H���:��wh�_�Gpm���t9^�t�d����2F����R�ؑ����Sk����B�.�R��r\�Zǁ�b5������Ű�{�lQ6�5���{^��y�y*�s�|u6D� �N)�w�����C�g��P/K�m���\�F5���A�?,j���A@��,Y�����gC��㛾���(�[pˊ<pq��r���7'�])&.��2ć~?���ϧ�Ї~��-b��g:%�������ï�:4֨	P�`���1^6�g�u�Ĵ�o�Jq�"�"���x�b(�$��<M���0�����z�bْ'U�p~>�f�����ӵ���H�W��
9ħ˱<Ļb`�$͋p�
5�AÂd]�9}V �Pn�Y���]@�D,}�.7��g<��e��u�ll��/)��/��z�JIj�>�c��d�`�\���]��^�EK��w$����<Y�ց>�Q#�2,^#����DK�x*�")NP?��꠱��j����gL��I�+�P|q,�R3�)�/;���FVG���	i���y�h2��Zxxy������.��u�X9�i��X���ˈB�[�K�Tn�4/
ٔ������"ۊ��ꛨ��?��:�^-�X�`.�i{UZa�;���k�5n�)f��BL���ުl�?d�����ޤ`�X��:,��y�;�,�Ђ�#$�TEb枂(��5��sC�W�
T>c��X�C���;�����U88a�Md�V��n��T8��z[��Ox@�)�o�z�]yQI�����9�5��?�g��z��$��'Ǥii�7y��#��"K_&w3��W�W�c]�'eL�{��Re��@;�`��۩g����:06m�rc��n�P�v�,�������*�`��I7M���ƢCj]̰岙$J2�N)h�q^��{��+~��Ջ\��t�4 a��(ǕL�8���g��6� s���3�,����?��2@�t>#�yMFxMZB7�̲�Э��K�_naA9L�r���a���:����U���)���bi�CHkN�S�R����Q�yf�%-�&�O�� �$���6V�L��  ���Y����|��E��F�p���x��X�~�?�,��d�x1�넞�����A�1u��"��#%*�ч�C'9y��d�AW�8���F+Ė�	��YR�J��=���i0��[��^4�kGwZ=�3i�Q\�>�&�0�)��f�SEH����<�N~��Ը�z��%���[a0n�K��� ;�`��o��Y��BI��#�����P�i$hOo���m�Z��1V���1���ɷ��6t��(sv���X-חt�]a��]��?4��!���ـ�n�c�� ЈԸXlxVHYEB    fa00    1e20�8i<��F[��:���)�jҿh���yz��b��=1J�T��c��w=@������I3F����T���-���=�������q��T���)>�z�U\;�q�"0�>;�M�Im̯
��lP�8�̺_��J;�e��wLr	�f������p|K���dF]��7��dt
��k��gT�VEb��I�$�1?x�[�D���F#1H�!k�������/��7��8>J�1'���z��0�k����@�|��#(�0$'�;�e�rݫ��J䕐����^}���jWR���Kë<���}��M�);�^�ٴ%mձ�ɍ�����WÍ>2��Ж����g�A�����-����K��H��xLg"�B�]d$J�$L��Cc��ꂾ����ݟ���'$��Ե2�ܬ:�'���8���
�,��yf�7����t�|�!I��+��8^h���H����v������_�V��x�8g)�d~�[�E��q��BŢ���~�Z��\�*զ��h~��ag�����;xv[aM%��zq�a��L�����4l6�24�6j����'1�׏Ն,��J"3�6��
��'���	F!�Nu14p�a�r��0�4��Π^�`���u�k��:l�-΅q>��-2P'��r	�7��r�R��h����0� YY�~!�1�NB]��0IS����F��-�2ݱ�`vC�T��y�[�.�fGߖy�N{�hb��=p�ap%�Z��&���U^Gk#�x�.�7�����
*E� OT�IF>�}��K�C��&A6��:F�V��A�F�碨w4SP#��(��s7V�҆�b�B��ԨV/��&�2դ!�����F�5Rf!�"��v�<��:��U�s��ѱ/��S���m�+E�d�]@aU�nk����3�?�7։N���5�"���,W/m��]�~���������g��ί�7�8�������#�}ex�΋���['s������9d�m�9��6��,I���d��ޭwXq����1�uvw��yA5��@&l�˛�oA��oA�z������A��)0�=�S[�f��w�gThw��+c:&6��*M�8��@��b�������Rqn�!n91.�e���Wy��8U�FҀ�"�_�@�h�w��y�Ug�?a�m'� �!��{��CqZoGƋ��J��"��P�FTx.?SD�K.4=�B=�K�%��X�]q����*6���'Bv�7�x2���1)��=w����>XN#�c_�> �Ji������ˇ�@��
ĆO���%���r��y�L_��Pm9�ަ�Z��$�| BO������� ��_2!����0/�(X�~��a9o�*gNz�JVU��):�|���ˎ��i�Bǿw��m>\P��ۻF�!��#{a}��d�}�Ch��]=W�d�ioWa��n12T���b�ʏ�7�kX�G�n��W��f�~Nۊ¯�Ow�|�%N��ȎEFZe�L��u>�O�^����E+
��r���X��13�z���	� �t0�D�(^��emH�Z8Р��Lxz���ܗ�0�U43X���)��)b��4j�5�,��,"I��$j�FN�+���b�6f0��F�]��)pJ���i������m������'���͖�Z�ė�X�fA>�o�}�4y�T�T�hv����p�w�I�����l�7<�)��� /e���+�˾OJ�e|���[��<��p��1e]�G�D!V8�i���ՏMI����9�͜�!0�����^�Ʌ�����P`�@ȭi�Nq����ڃ=�!��:Q�0U������+or�<�-�"�G[p�s�	~�"�SJ����^j�DT�� �^�"[�>�dݽ��lܲ����Y�j�����3�:HA1g��ow�|�C�	�>����,����/�1	!������?m�.�`�1p ��k��د6}��$��`E4;��[�,T��q�X'2W�/��TN��2�A>���f/��R4����n��z�M�x��e�=\-0o�/��=Ӏz�J.��I���a�6�@Q�(�ԇ,���0'4����q������;���3�h�-�u3�yˤ/�^A�_�A�?d:Py�~��cM'��pT)��6b��f�&�S�t�/ oo��tJ����S�(5̏h�;ͯ'�5��O��h�����\y���@H��ll-�x4pR1e;[)���mt$tZOi�Ѿ�Z3�6���)�)��t�B�����4���B�Q����]Sy%�Z��h$Dn}nN��	)>��T1���ܛ �[��~�g���7?�82X#�;�FW[�4�T��6h�P< �0p�VC['�v.#�F*�K(�嫤,��ŬƵ��٠��RO�|>~�9h�> V�Iaد�#��y��x �L�8d��=�5'�4�E �c��jy�����U�*CC��7�v	mn������S�:$�nh���]2`"T-2B/ >-]�oi�"��^:�a���k]���;]T����)]~/a�4���^O�:����hd�֑��<!�ΪU?N�(�g�HCv6������O��یS{�s�B#؈���|���2��o�&z����	L
�&��j��L��������[R�,�ߢ�|'���7���Y�vh_k^�*X�m!g/-q�D��˥�&\쁀}��V;�-A2�����҄�.���|���/1;����Jf䂯�5!$��b�60�~����.X����3�Wh��t5WO�+�5�'�GUK��c��1֩FY�Ųxz�eÆ��X�<[sa�7��޷�5�90Ԯ���-����F�FZ�չ�_�����X��6r���b�r��&<�^�Q Ka��^�ys����bOĵ��D˭�[��/i��n��v$0e���,J@�Rge?`@�]�zm1��lm��	)�1�ɝ��(�|�n�;<���sh����L�a��~(�L2e&�}��c�^��t@�1���i�������v�R�ec�@B\�g�(�����:�3��<e�E�k�Q�����0�>�UԭI�XC�xg;* ݠ 2�M�v:F}=璜��E���f�/G�.:��6[�l���:��)E��׿j�0ǳ+�$�28A�A7Ύ)�f�F���A�Kg4j��up��_Aɉ�ۥ+4uh�pbV��C�C�W`���#���u$�ɞq��M���_8:md��jx` �͇�'�<�1��}k=Unr콭�V�wR�0�l��[�a$�����[����ʅv�/#�S�X.��MT�<��Ĩ�����O�)6BQѸ�A��,�2�g�H�q#��h7u�d~����	����c�F�����a�.^}�X��*z���zl� �S�;��F���|�?X<P�^C��Β�v'Y:%�D7 hӌ.�����?�׬?�}�`��"#��j���` :�n�eo��hjU_M\Be�;W��"ՍB���n�Xi����.�&+E�Q��[9^��P�����V}O�\���8){I��W�#����V��|t�Aѳ1��~�%�-j�҆�>��z�/f/��Uഔ�F���(�E�ו�^xP�\�`Ђ���+ޏ�dhxqa'�p�^fU������S� eϩ��G\�/����+7��k�/h�a;K�>��Y��e�RoU���&o0ѡ�ol����bV�q��s34�Ns��?B�rƗ��/��tq�
]Ƴ\*A��(��f{�#sQ��l�5J�5Y.��}��(E�e��u�o�:$:���䇎��#�"ha4�T�f�j����	�i� I6!�8E�9��-HIf(��U�쀸>�.ҝ��m�C�F���|aOA^���K�)r�UUmiɤLva,I9�<�P����l{��(����^�E���|@f�Ω�����UW��������K@~��{�U�+\�=m��لlң���U�Jl��n�zZ�c6r��vU��p+[�"�o/I��<{�Q8��vB���&�5��g�!�}��V���Ć}�zH����E�%!�,��R8@��6�ۂ�_��5�:�y�a�)uL�ʡ�e��fz��-�l�C��~��A�0��j�����0_}n��eUC���r9��=�5rY3���T�V2m?�G���0\;>��rf�]GFKn��	.��,4����v��72�#��A!kg��.yND!S3�����	�c���!�1�s9���H��$[�	:V�=��3�g�n2�������j�$����}��9���E��Z�G@�ʊb��7��J��}���I�Ⓢ��9�9�5s��~��`�eI~�����צm�%�E&�{�EIOmMGL�L�D#�r_�S GFg-��/F�?��R��k�8�I=:7��h�!��N.�p���I�	��6�U����.x"�f����5io��N|��w�Y'��Q� �[�x�_q�?_z_��m��x�z�ӿ���Tκ�W��H��3=x���qdۆ�y�a�Ճb�!U��[����@-����L]]�dq�1�s%�?l ��dA"a��wML�ȼ�x?Ӝ�<fH����ȯp?���|��ӄ"s,����Ș�O�
�����k?���_��J�2MZu�z�<u�oFR��F���d��;�ɢ�rzǖ�52��9,g�5�x0	��� ��O�x\�]�.�>�[^�ڦ�U�^&�f�5�O���J�/q;Iz|L�'J���_���>\Wl�_7� o���>��p_��Y���mg_˓YC�&�{�1�l�*l��>��
�6�78���|�!�m,!LL��;�/��s��уCX'Lx�x�z��g�
^l��.t��U �Ю����n�w gf/o��Q��� ��l#e/)��8ఴ��Y�-��#��X��;F�
��)��mGZ������"w����M����.&H��Xܢ������Roz5��k���j|�f���g�Y-Z��A!��QS3�xs+����1 �Us����ǆx��4�=yj�o
��#�ev9��Sˮ!�֨)T/]4F�1�$��*�	�4��%�P��s�n��7z�����;3q��"OR%���Qo�� �Jw�ۼ�t���Z�i��ҕQ%�F.��ơ��G��=|�m2�L�mH1�y&�1�=��0����X��bN�w�k���0�1Q���
A�Ůp]K;���[��̘�&!*�и����脲L>tE^���ּ>��m��Q C��4	|:;b�h�M0 ~�i�����(�;)�Eơ4�woqg����J��Br�?;N���F��Z�itTv�y���h����Rh}�ѝ��v2%4`j$GE�[���t怸����!���aÂ�fʻdr����7nEv�8������H��?c��b��0��2��1I)"��f"�B"�Ќ[b�G�>@vrEX�Z]���oP�/�.��||���x��M�TT�'��w����n
��1?��%��0����e+z�*�X�ݤ��'����;�C�`�Ew]k~���g���擄߸oo�L�{ZR��a"3�/�ˮ_8^��b8雎6�xE��.�#h𣯵���.�'���Q������\���Uy�����p��Ω����9������L��ؠ�Hj��q�J4Wy=�O���B�p�j�#�����Gd`i�z2Y��ő��P���ūf�We����+H�!�e�b@e��1}�*����3�KQ.��A	3�L��R �:�����}�D۲YZ��F+�Cm̴z�F)"Aˊ��2WkI-N38A�Y}� 6�쟩*�1����%*!�z��d�����ֿv~j
���uL!��-�A̯��ꆧ}��l���@bM��O�)7&�O�s�P�o`�-'��W!F��$d���#�~�ѹ�L�j7�'�R�����a��7n֗1٩R���8[���s �&5��$</�b�.G�ku�m��n�,C9�S�=�	�-���D=����{����q�w�/=�X�\vE�=N�b,4q�R3?��s��tCd�+�WG3��^�u!L�2<��W��-�Z��i�k.!۳�шCU%m�+ҨA�/�Uv^i��
z ����Y.�ˡ�&2�E��}�4�]nh�:���>�_4GQ���U�E&\�i��B�!.NP���"#���a�T�Z�I��Iҟ�`��="s:�6�G�n��g;r����W��R�6j0���|���ݚ�����0C3�J`̀��_�pC���	j�1/��������;���ht�Em$�a4s/�����I�����E@��_�����?|E��r�kv6V�z�"���ٖ8�T��`�RE�yGIg&8 ��|d�<�^���U���s��5��ȵ�2<�j(�h�B�B��}.��!Q�@Xzs�"�C�����	l�F��^VīlL �Z��f��r@�����[W�"nn�-�"��Q�,9(o[�T�&	&�lp4-&��� �	���[�Gt�3��]�	�i��Q2�W�*d7"38�
�q~��'�ݱf�5�K��<ݽܮ a�,{#�9�Xt*=�aQ�a�9һW��%�X2�A�|�hbF�+�+y�J}a�_!�E=,j�ޮۢR���b~ˠx�� Z9p:
����'.�������	����vb��n��N�2�U���S�7F&����`��g���c�-{�ET�b	�����x�8�y\Ү��DX�����׼�$�}�����l���փY�qwE����M�\"�����B����E
��T�X�u�X4��E��-����<O��' ���R�3�^,JY'�Sl_G�K���H!FW$���N�;~�4��	�t+�E�g���j��f�!�9���_��1r�[������G�q�_}�|e���n�P2@.%��#�����v��S��x�
p������C��3�ay��M��м�4��o˫/$�'��G�����r"�EL��%bR�+�I*E(��S��7q)[�QѬ��؄�%���p��u��n��A�5�=��<�H[u�3�[^¥*[��>���.ҫ0��k9k�H�;n�2X;cj���m�j��5�4�����D�Vل{��N��_�������+�q��y�c��P�d�E��%���K�b�k�3���`�pk�]����MA@� � �G��γ���oK�;�����t��w~U��ȗ�j�U`&��$n_��l1߻�����q���t����M��]RQ�&O�S<mH,�BF��ʶ�[�C��X�#V�[��z�R+�Y���;�&��ͳ�p�~�ŗ�շ[�_?aO�L���N�FP��ů�@x2,)�&�"4�UYH����o|���" d�7m�Y��b��N��a�x3���=@�^=n��>a��3"�G�~�rf�NP�k<۫��&�H�KAA�C��p����ZV�R�Ծ�⇳g�ь^��Wf`��HfvRI�2����[ �4��N./����"�������幊,���yM���
����~(������{����A��	7�FXlxVHYEB    fa00    1e50�b�Bt�`E��ϫm���A�w2�R�JA�ⱃda&2Xs�����(.�3��o��!�������c`�u��&��Xl���a1��9�����.6�
�e�"XS�$�W��
H/�Ⱥ�2IeӅ��k�{Ͽ�re��^{��P��#�&Q4�^t�,Q�)��^��$ ���lu�$�p�x*�s�|;ۦSt� lOlZri ��;��������НϺM�-�x��m�|oOsu��_��ZyQ�j�eȮ�Eq�˦P5�����A�xq�,>��\M� �|^<�S;ׯ��)h���2T�����57�8�O H%΍����g���/�>�J�G�j�`[IX��}�R�|�Or���ROs_���}�ee9gs����������Ad��Ck�;}���שx�<Z�������]�0��U��3P�%�d#��)���ܫ�@�l�[��*�	�T�P���M��vހm����Y�[��t;h��%�Q��cO�εD����T�o�Uv�+�23EB��9���]2�֧w:P��A@b �� �� |�JN�����<��.�`Q�ѽ�,��J!]�]Q� t�}(��<�ϫ���~��}�q���ٹ3�	$�28/��7V���V{7F�FU����W����M�;Q39k���a��y�H�IlA|F`l���˓��?��OV��ï�~�\0����Y_Dmds�E*�8О� :Q�?Pp�����_�i��c�����X^U�Oݣg�i�����q���1��HJ @M���k�	L��wF������"9��3��Z�����\��ã���Ŏd��Z.名-0�rf?�#UJ��_�����IFA�|G�T�q��RD�i_�f��3P� ]A�.��Y�,�O[5T��`��{�*)��a^,�=Tm$w����V���rۤEb%V^�Z-�<�&Th���&�s�l��l÷|d��0��ߦ 2?�V�8��V^���׊@g�y��L�o	��P{�F�|�eH��؛�ݿ���?�8r<0?T���i����$����3�Q.Bȳ��-z����^ě\����I{�x��o����m˴�;)�)�#q�z�����[�u!9�)�6�xi_�l Z|��n��2`v�{gD���̵���H5���
��jZ��\R����9R��h���v�r[���0�F#��9��(%�th��/��R��\�a1#���m��
�5jD���7���\��.E2a�BPS�
=�W%}�|�S�IT�O��!���Y#�Jo�*�v��. �_�{ a�7�U�ĆNۛ3���ܳ%$n�wy�"r�%~B�,��o]g�x2Y����}%#dm&�8�0Lb�ˎbbR1��)ܲ �eU�5������n��;lGT �K�"!��r��ac��C3�8��-C���b؛���~[Z	�A�{��x���#E�'j�`�Q�D\L$���g�7�%N���P%Jx�@��E�H����<	�8�x8y�r���L����m�h��F��>^���U0'�������u�사!�N /�}Wh�J�@7��PΕ�-�� �KG�p�&�Q���j�|@�t4w��I�И�.���ۈI����3 5��aC��N��5&i�_�=Lg3�"�:����>��ͤ=���us��Q�Y7��/���&����X��?*���ty�����[��XX��G�$�G�������ua�oM-L禵{�Ku�קeE���M&J�� ��8�@���(�T?r=UC����I��ӟ,� o���W.~����'	��j\����%#i�uk�x�O�\h޼�� �I�/9d�~?VFx��Bgda�G�ɕ �T���`Qib���������-����L����y��x Y��s�[�q ۡ�[�T!fa�o"��{��\��@3�.+��佨��g66����j\����L��>�oR�R���31`<��Q�3�R\�}����ʢ����K7�� �>1!��k����!�~e�)f"�e��j �yK�#Y���g�5��6M�����UT)x�9�LB�3�Z!�=л��>�E��y��&��]��f�G���4.��1��
��g�cT�̈�K�}�9��8�V�:`���r9��: K�L8!aT�?����p�l����\z�8��O~���1�M@��A��)S�7t�E�9���/���V���+�J���)�i;��(	ͨ(��iۥ1룏j�M�w����7�[%���I.0��C�,���0�=�/�ކ>��3�$
�������F�=���Jz�
���y���p�1l��aʁr:�(> ���ܪ���jۺ#k��)�gz����L��5=�)����=��� ���b�K�[�/�����J���ɾC���Җp��[r�ԑ"��y�5��9*n�A�R��
{��,�D���"}�5%�09���~��� ������~�Q4Wr�zF��rY��	_H��P�?hek�&L!�6�3X"��jJ�sW�����'^�^���%��lQA=G�]���}m��RW[Z!"�e�`2���4�����;h��'�A�KI+Jb�vZ�S���O���+����y1�1��x�ź�����B���4z���U��(�6��je�|Y��[��v���Z�;�,�+����e�� ��Y��D�_����d)���#`K�(����O��Yи��hr�ד����EoϐEl�aM.W�g�u������-�k��o�~;�}��O�KP��j�\�+��8k�C����%�Ąl�����3/a��k��~ADQ[H߬�
�<�R��L����#�s�qD�yCl2\2*-<d�ft�I��=��t�9#5j*sg�Hk��Fbw�J`R�1h�G5t��)m�3o�Y��|���xD@���I�5J��~a�M��i���ɥ�Z�� �0�������=a�����]wF��~+>Xs12	`��>����Ѫ��������TI!��fV���G���B \�"?$A0$����AC�xː�A����}�g6��Uz���������7*#DP�e7@��*E2�n�%<q���٣Y���&oS
$)� �B�I5=�#9?X��a;�X���Ҡ�a�q5���?�f�vA�u�1�/sG`|"Y�Ϗ���PG��n��E&F���՚�}���_jZ��`$���-Lݤ�������^�C�Z���Xa�m('�觎V�����+���l�U� �X�6ߊ�B��W^�I�׵����}^5��Kq���i[��l�c�AHU��{<�X;2��f��	]3P�#�La���W�WB97�5|\z���N���Wh��1@8Ӯ�B�<ȳW�:i�=�+���ŉg¥XA��1���76���FZe�k����2�Kotm;	CV�f27�C�	���љ��7���Β�K�f�µ"�$�B�R��[/d��V�	[J�
N�*�X�Ct��l~-1�z]��/iws�?�N͊q�Ӵ�cٔ1����u�,��7&SK���ٗ��blݸ�|�L+���b�1����Q"=�^b2��'�~�ie�<&?%�v�)�:�m���J��<�Q*�p���ّ����JIw�_����Z��!H�`��K�����Z@������G\�[���ݤ��iU�/�M�����d�W����Xt�P����:h���=?`r�P1��|g_bM\����du�n���9������s��{��CJVi�����j�Q!t� Q�m�J��ݚ�7NجV
��R��)n�����D�#�㾝mp�_X`z5���>s���0/|[�y�?�$��aD�5,�UJ?���]֠��pǓD��,��B�/PT�r69E'C�l�|�l��J�t�.HJ�g�{j6֤
 (N�#4<5S2Ǵ�}׼���3�"�I�rP�/c����	��p-z�A[9a/;yTO�m�K-���;#��� ?�L(|�mg�R8��O������j-XcV�ѝ��-B�����T����KT	�����_]si7�RqY`���`�@C�vGXiǳHٔ1A�|-֍�A�A�Y��뻌շ��Aiť��!�_!�����t%ixw!�	^7�.ÙNTE��C�(�u �G�hs�����:�0mX �Pz֌�����c�����3�Q�i��y�N�p�Au��%�I�"�˪}W�q`�����!eZ=
(+��.��YH
�_hU���V?\K����$x����d��:�9'5�,�}���s,mQO8�;���i5����)Y����>����V)4W�=��j 0,�)�����]7ֱ��ʤ�[�v&�V��k�����.�'Y:�ڰ��¼z�{�+�ҷ�+ĭz,�4t&r�����an�l���o2���L���$�.#*T>*I�?��49����goBG��ר�!c��/&z��@ӈ��P"�����4�Y��{qW���|h�0�D�7���H�"��;���^�p��2��j�:w?�9c�[͡>�r� E�/͡}� .��< 
��B��)8J�Dc_�:U�D�c���br��񈲷�rJvV�P0��߽GJb(�h9�ɕb8�N���QP����&$M�K�{��� cG��Ϩ�=��W�,+�p;����]Ԏ
��@�{�������lʟa���Y�Z�l2Kf�<y{���r�PG�����y�Yp�Z��~�1�B��r�ӎ�@
�C�_���� 1�JI�����.�Z<��T{��U�|�4��cX1u��:nZ�Z��O��k��F5|�`iѼ�]F!��o�V�����$rUp�b�W7��*T0v}��{���UVUo���Y�r}�p�|�y�kf��N�<���̥�HC� !�UT�B[�=�ʤ�+=���j�V]$E��"@�XA��֔���x���r���i�4X�n����Y�9;=_�4�\i ��#�Ǵ>�z����~K�Y���Lf����A����5�aǺ5,4s��Ņ�r�#U'KϦ *]��P?�e{�芴�ʆ�#ܖD,PRo�y!D�/��ٛ�l/��c�H����-V�5������3�r��	���N�.W�?�7�����6��Kś�,���CO^R?����w��_�K�ȑ�X�UjDN&W��\�0�����- �_ֻBJ�qS�ݚ�;�sN�g!s$�yf���\�	F}o�=���j1�J���f�Qq�����i�/���
GM0��? �κ���>�n��aO��D��$����?����_>�^7����#o)2�ўo�k3.�����1�n�9����}?�D� [Q�o\9J�4�8K�Qo���:���שּׂ!_(e^���	�
���{h�+_�~�X.�@[�$���|��g�&�U����:Te�l~?K5�<c	%߶����`����wm�rg��$$��.�S�賗zҼ�5�p�pG��u�~ŵ`Ζ��}ӗ��6{�|��lx%;����s�k�kֱ�fNo�E�'�x>'�p��!k�Gg�O�����"�\0��E
ω�:����CL�hK
B${�����>�uYY�e��T��5�۩M�v�"�]�C!ܭ9__P3�\	�ȇ��7\�ܫ��Hv�mw]��:�������C���7{�Jr���'Gzx���=f��%���7���PX�aR�S�|�_�����q�����Z��-���N���B�fs�c��{X�'J'�x�<�a���G��k^�>���˿���bZ�<�y��v�6e1�Yy����������/�7G�x�4��%)��ͣ�/y>E2�2��!c���"C:.|�O���kE��9�JL�����䝒 �d�R�;o�c^T����7vt�,��ޥ˵��/ j���"ַ��4o.iK�ou�r�OV���hUGk����1i`V��I�S�J���ն��A��0��-��k��1`�6����K1&�C��0cӾ`O�'�����_y�`[�T;7��@�mZ��(n��!*vβ� *Χ�%4v!���utw�ڰ~�c�x#c��N��&ʚ��+ۇ���@��� �d���$�N��4�X�5\yFp��c���FջQZu�����L���h��]m��@����`�O�S"��(w��̈́y��$h|�W����>�&�|z����$�7Cn�)�-}�U����8��|�Ѓ+'�䃢��/<ʹM�@��۷}���#���a���I�ir{�+?k*��w2?�V#�b!O�&A���'�Y�HT,�&�����M�A�����>8X����hM����O:��6T62lSw/���o��ľE��N�B��{�щt��G6W`a�s<}����ɗϙ"�)����ħ�9d`Ĺ&0�D��μ,�;����7�6l���q�=QC����ے�up2%WP�j����E��^w�.(������~���BۄK�C{.��d�!������md��)o��������D� �E@mHm�m���?���.yd�s+C8��Ǻ""�{F)�`�B�8)��Ş!����ܨ�5%c�"O�(Up#����<�z��w�^X��S��
�PG�}��F/��c�Im��>
��a�ݒ9e�NQZ�r@c�?��ީ��d�Xٷ�DD'�	�>��i���eEP�+ w��91�pݏ<�#�p���m�o#���sE2u�u�!��5��tRP�D>� -1�K��,N��ql�7�1o�{�!ma���nkIN[��� �_�X?)
��j[��Ϡ����*� �Ȣ�cS%����@|t������ \x?��%Q�f��P�3�Yu����p:g:]���ވt�3TG��B��v��������n�'L����c2ի�����5���������h����sW��9�<�_$��B_��{����i��}������w C�/.�b�N�FO�'&�l\;]H���p�h�n��DCRދ��t��F��烳���H�e��H�bK@r�52\Yh����)����$~q�I�LSJ�PC�Mv\T�����#:;WWyo�d����DJ�=��8ZR�0\�ט,zd}�d���F���ҳRh5V�xP+?O=��Z���T�[q��S���O��pte����N���[>�[�J�z�FԺk�ho��L���-j3��A��b�d��n	�����oC��4���C�F�e���Z�#����y�uJ�C&jH=#��E��En�g�4ص� /lfW�3��;���nY��U��ɾ�p�L�Y���D�^�Z�PH��1ثJ�n
��HXo8����DÇ�񼏓�*��^���_����y8���!� ��d �NSKHJk�4��@����_|�W�Ɲ�߄���:���U}?Uj�%�������*�zV��):Rӡy��"�j{u�V,.�V�Ɵ�E�v�GDܹ&�h���[|�bi��Z���pQ=��Q���y����#�ө�%{����+����x�b��,W�,��M���>�
ӻ��:��b���n^�I�IN��3��Z8�S���DQ V�R7-��XlxVHYEB    fa00    1da0�sε�L�����ɧ�U*uݖ�YV;jpd��!%�+�z�[q��jӼ��Mw�)���v���@�B}�&���4!��W\Z�;ʭ��)`�,C{ɬ���pd�^T��P�Is4������6,�^[K��G1֕�/��ɻ�q�\lc����F4J
>,��?�7��29���Ѫ�k}w\���?q��;�)�=�t��w3��Zp�\)�\�
.��%f�zu�WZ"��p��!{h�K���OM��w��^&�����TƊN�p�ے��6t�lI%�%z32������"=fj���7D���n��%7��Ց��P{lW�-����#�fv5�RҳA�Zp�=��OTMQD����O�Q�
���A�Ո#�2�,�+�r�8B{$eEJ=�����ԽaDů��SK���g&|�iS
|���a8����s�q�r>�ۘ`I
��B�n�Hq`��+X�J�ʖ>�Q�������	X�P��K�xE���}�;"�k���A�Zه+0��f38����ǔ�Y9R W7���Y�~t^����e���
K��\*�
F�'׌�蕽��U��L\�l3����ܠ����O�ꠊ�ȯ�c�s>DI�!�]5u�uw�O
|�.�)��ᓮ!{_%Ѣm�3(��v~�b~�[\���Ao~;�3��޶���ܔ3��Y��	"r���n��T��|�g���%�+Di����N	UWB]���K��E�d����
<�M���&�J�dx��͇�~��9�.�h�2'Mm+�d��B�Z��st�6+��G�Ԫ{[����8@H�t��sX:7��yS��
xԛt���B(�P=��K͖�H��U��qu�XRÒ�	�>�
"�>���S{��#Aw���{,�n�%W2i��,��"�>h����+��v�:��X�:zr$I��b�{�M"�BAmW�7�=K>dQ-�BC�w~�E�"���e���F�����	}�^�ݣ�[�"�m�R��g^��$4���t�0D��
P���b�}`��n�	Q#�b9����m��B?��vlWZ�K�q��������	���Ң8�F5`�ƃ�o���(2��x�{�ҥ���&����	��,a߂c	�+Y3�
�+@Ҩ��i����	|u�E��wa�O��O����׿���i3�Е�^������5[����%���^!�i#SWIS��#��:Pc���c�����Ka�����*P��E�yq�λ_^�m��E�ܤ+K*XA_X	}(̓5�K\_'��S��EW����jm����jd��#�P���M��T�� i_����zi���K3i۲��Uw�]@�;�p�ƞ���1�S�ŰB}�c�Kb���μ�� #��[�%1��Ε���@Y�ξ~`���aw|v������u�ĠĜ ���|&��L�Fj���ς����f�YvT�@Sʫ��9N�6�B����47�P�z~������G���.���n+^\F�����b��ʳ#V�9�'��˕&���6�˶��ˁq�d�����p��8&��V�S��/��/���� ���C��$
�'~�kEQ�+eTͶk�wS\e�����X��{Sk��R�Q�,J$�t7�r�Ρ��x��z���<�l��ݦTa�"�� w���J{��^�$j	i;7�� őT�R-��ʵ�zPLi�5(����BT����`F1�e��l�9���P<����Z�#lS9;JI�21��9����Ϸ�y��Zӯ�u��Aq.�xN"IE��Ϻ�����k~�0�8 �gq膘z��4�_:dY+�	�DW��:��#�Bk7n��c1��O�B�9<90�b�����o�l�B�	FFp��Vs(���5�[=1d�QK!�4�'Y[���������ܴ�x�_���FQ�.\O)��<�z�i@��B2��~z��}e� p��K~�[�8�˿�*i�ȤT���~�䍅&M�?S+ȭ���N<h�R�N%�i�L�Qj�F�.��p#��w��0ʿO/N���{��ɂ�7�T���rF��m�fbY/F@��;��CtF��=�a;=���<Ϟ� a	��g�t܀�8����?�
�=�XVt���|e}a�|Ia�}g�8�s�nHBc���:$���ֹ��A���� �t�Fl�����5਩?��7���+�h��d�6S�+�
��F��$�^갣b�m��	?܄���zNU��B&E��yd��
q֋D����5�gړ�V%F�/�Ah<�x�k������s��)����Nct��?,?p8��� ӂ;~}�4��n bv�� D��7$�#������ ��cX�WYy�	��f�T�0�8�jy�����e6i�$�u�$B�x���E�Nɡ��@�d�j1CNqV���6�S$�=@懢^��l<sDWZ��s����ͳ��B�?	�����a+�E�T$1|-�����?��o�bo�B�##X$���DO �f�5}D<�0T��c!)�"���+/n�]�Ի�տ��@��=`�q���XK�i.��)�{_G���5�OKy�.�Z>.Yu)L�������PbB7f	r`�!M�UmAHW�*�t>l:��F�B��ι��Y,eQ�����~�y=��G�q�.���Ԅ?d�g��E��0�l�Zk2�PR~ !�F�V�qJ�`7u���������(�|q�]�M�zn�d>�����\��� ���4ᢋ�B����haQ
� e��2?.�zh��Y��/�O�$���am\
�7�+���F)�:����^V%<���P]f�4m���;K�<G��Y�������\z�m�c(!w}�
ZK3�wԹ
 ܌�i���'	�m���ed��]�U��ok��9!1[P��A�����DD�WsOa�]Ǵ����]�v���N�U�bϣX+�ri������l4|d���'+�y�۶��Z�[�x!(1��N�ƀ��De��_�ud8ϔ�݂��=�	An;~\�N���E�X]\q���_���o����{k��Y�Z�4Qh�tkEW�ز�e���4��Yh&��`�o�}�=�_�6����;_��O�T%$*n�֔�1&�Ww��"����y��p�@�R�ǐ��H%���Y:9�6�����!gu��6�/�ͳ�=ǀ�����%s�[)��s���D��@54u��[�d��:Ȏ̼�5�����g�S<��-�8��E1a '�`c\�1V����-\���f��w�QV�>�hT����f��z�PF-yY
�j�,-���]���ױ���$�m�E��6�e:Bk��V���Y4��,6QQ���f_e�����!�	��p�iF��3��sU��>c���-�3�'�]��q�w�aQk��^~~؞g��<���4(N��e��V�:�ߑ;�h����ͺ)�d�[2!?t/ "��G"T�W�w
��>�d�L��-hgs�����ӊ��tr��|��'%.4�b[�'Bt-Q\h�@.+N��~��D>��^��'�꾃�P��
^-q��We=�vð�1���kQ�h�D
�"=�rc�]���E֌��� �mn��K�V�QNP�m�ui�d�Auƍw�P��h,غ('��yK�43C�=} ���b�5��
��U�����X��ǩ�2�Q0��J%�1�D�[yq�9����3@����tR��A�
6�\rw� �2el'vn��15�Fu�EW'��Xր�J��<��,�HT\��l�m9��a~����iM�n�[{�zT0ūp��D�V�~��@��h��KK��Ԙ��Tΐ��)oZ�ƥ	-{ǣn�%��� ��AK����(���u���H8,f��c�O��ס"����Rk�Cʱ; ұ�fP��0�Q�>W��2#C]���8�8`D{�&�ub�ӄ?'r;���u��Cg׾Sic7P(�5���'�ۋ�n�)V(��\�[��f�~�Rh�`L�+T��sѢ�
��B
�����f�TP{@)� �Л"�Pw��>���*���@;�F��<�Ӆ�Gz��@)c�۾�^|@7��=��D�~$,�f���kQz���*��� P��[�6��ԙʸ���)]�<iz2wߝ�qz��.�g�B=�
r�?C,��_��$�"/k3�t�8�,�}}(͌P�#�I=A��"�)��#\����[]^BR�x9J��5_���M�B*���1�h>,�R�|%��#��3�j�N㟿�7^�NY����rg~��7Q�"m��Z����'��-�U�G$���<"���v�(�۪��/>Wo���jK�m��sd�	a���=3��t"�;й��u�g/�%Ջ�ܒ;�Z�
��^Gr^�nB綝�6�7����� �}͖w���ثݟj��ro�͓�\����BU����ܧ��w&�<$����mN�gYC�9��vӞ��.�M�f3n��T��Px��f��B*B��bVp��H�xFuC'��H��9.Uv-.�-�񒺱T;p$���`���D}0C�M�x�\#��荦y�N ��-tx����H�H5�>*���[��|gb��O�^��d����Y�Mʿ�� ������˥�~�\V{s�����,����zS���v��g0�搨�V�v�M14�-(
b$�H�V��Y��X_t^�Ԯ\i�I�\D���Q�빊������q�������<I� �ɪ�d.ݵ��ة�hjdD0��?61�=aꡠ3y�����ԣ�M'�(p�X������G3ͳ>���-KP���Ӳ��ˠ�������JC����,X&�!w�Vo`��[�4K��]��w��k�<k��.���ڕ�#�y��-MyKe�N��<d
j,5O֊D�
�;���iۅ������[�y��'x��J�^���"X�[1$�X!f�idD��>�T�c1?a91�0�����Z`�e����~ү���dj8���i�<�f�r��$#s����v	S�-'l�
����|=AiQm�Q��22ַ�Y1��A�
�E~G\���)}\�!�jBC7��:5��D"�v�
J��>�׍��RՎ�A��^��&Z����� q�t�ftA�P�v��-<k1-��l75���D�C�L"�qD����<Fc�8���/�y���[�\^�k�Q�+<_>F���')��	��jwx�>�����?��`9�rϴ�p��Q�Y='!2��`������}�<��ʥtP�W0��q.�� :�Lfp���?$�d��P _��
&@#���A��pi���{o�6�oƶV44� lr3��Q}!u;��G�B�}3Rї�����fod�./--��f��D�2<?����Fd!|@?3���MP��Vȸ#�P9>�V`{&6&�2:���Eu����`yÚ��y�*�$c�>	�ƌX|�ҒxC�����T�n��}����r�*-rfw�^#��X�ϯ{�lk�ߺ:�M��
&E�g����u��V��x����c�y&t���$	���HnUtZE��xa߹!o)��	���哃��������La<H�-M��]���_��=��U������,��ӹ͢�_b�E���8��"b^�'{�@
�Dr7�X�VOp��x�z�0��k5�T>o�7�	��X��w��%Qy���������E�w��ls	�Mv�Lz�icTwG��9�`>�Gz���T� #SPԛ.J�7�w	}����TP�?B�}W�@�U.~����]�~���&��ˇy�M\������q����N�Y.8�x�{���)(h��~<w9��K�XE ~ʉ��Ǥ���Ye�M )3hj;vޅh�Qb����O>��g�r� �B�l>d�J�i\���< ���)e"rҰ�,�"��L��{V۫��gv������a�#��>p��A��>��݅M�8��I8sR����-����]�eH�n�'Nm��GS]�oO��f��[y������-*_��󥭾A{���∨����B�A�;�
�kJ��8qO�l�֒e�1�G��u���$�}+�T�C�ؼ2�=��y
��Npry�&�"��"Qh�C���� �5�A}��D���g���L�d�l�W��=��_�����?��JNZ�3��4@m�HqlIZI�:�G�U�@�^��Y׽E��¸���Z/g�|�wI��u+W���řnɅri��=�إ���i�I���v�:�&��Zi��^|��A|8��.{�tm���W?� �bբ�c�5��g��m�/�q���,8��]>�u'�?u������= Q�TQh�G����V�[`ck�zwy�IZf���A�JZr ���<dIq��[̬X�<-� ���Ԫ�W�k��PFx�c����B=m��7���h@֣D�Y�L��۾�//U";�!\��#&��3�5��yvmT����U�D�Eq�,i��K��&��+��۠���Bֹ�s���š]�4���r�WV�0���p��LC�)-�s�	�:��,��?��Es��6W�� �H rkh���Cd��b=~3�����̡�h�=`�I��V�%N`A���h��Bp,�^�ׄ)d4��(�CD���rx�*.����#�>�0ƦL��j"�\.+W��)��E�?���&�5lש0GӨ����x�N?����J�r�ɌyQ���#�{1�U�#��E���ƘcW.�H�'����.�7�7b,E�ga^A�Sp��D�0��A_g�XA�rL/����H�⛆�5�Uv >kY#G���m�^�OK�3,��|�	$�J=�Z:]g�v�̹�������<�q�:Xc�
\�3 �j�����bIb>�(��!�۰�@�`�5�o-��	���B�ѷ�d��n��Y���e��?���s�,���ܱ&�֦!���)�4�!_zӹ�mۧUkj��?oZ����4]5�_j
n�����"�˶���?�dà������sȡ8T<�������pP��ا(��8���]��n���{���	��-o
>�_1bH[X�k? u������"�":��x���.m��Oы���B��w��p��2�R@A���5���g��R�xA���nG��A����� �=- ���Zj-a�Tz����%X`8�7z��(c�L�@5�-䒌�Qa%������1!�"?�\���圿Z�-t�X0����7Z�6}�*z�VsAKI.����UBpN;]�����V%\��(�i^��B�ܙ������· ��5�h��0A�	�?M��sB���+9�Z�7w��X�׻���1�m�J��es�q�*�o���'�P�^	���U�HH�nl��&�x��f	� ��_f��`��Jl�
L���+x�yȰ�J�~���f{���Kw�rs�^aW�����` �+�-S��L(z2��נ�H�&�۽�cV�MXlxVHYEB    f314    1b50 :?���������U�	&k� ����(YQ�����Y���(:���s���$<0e'��S(򸒕[�Cn��
u����X�}ȕ�	�R6���H�x)�N͇c��6����*��f�h��N��Y�sg;v��d�� �O�>��n�E��Z̨ʋ �}<i>M����wo&g�z��}k�!8y����T#��hO���$Rn����B�O؂����)�5g�F�m��*��x������fJ+m���>�{ӫ���c���<um.��N)����_�/`��,z�ԣ�i���|����~���wZ�.J��up����������ջ�KyO��{(5#p��n�D���r��S���0-i�5An���GŚ�߾g��������Gr���!p>Bb���^�,?�oH�1�ԩ2q�����k�5�D�I(�d$1i+�A��8eI3kK4�v���B����n�z;Q�*T[�b+5�LX��#���FQ���:T��w��Y|���.T&#f�S�����d�C�{,�����e<ɴC2��E��K�P��Q�σ+;�w��R
"[����K�K-��9��T�n�����}�'�Fk��q$T�$�oy-�s�Y]��3'�KH�*��̪��p9$�n��|K��!��VL�4���,<���K�����,�N�[���C,�ס�Pg,Up��(���.�m��]�:�@��6��-��I�Xf�@)�->Z�pݐY1&-v9Y���_�|�ǀjkI��aѐ�����,�%hH���� �/B^�6uK�� ��C�������1.V�1��.V�v/���v}j�.��I��e��Jw\SK���Q�_x����u��*S��Cb�EȕR9�9��ڶ*�r�gU���&�,>����m��	K�2J1��$hO$,�o��x�[Ut~����k��o-WO ���2!b��-v'L��(�"҉���5�/������^���J�G�c�9��`�d�v���nP�,��{jb"I��6����B�Զ�¯��Q?��4�k��4�E�X�5�(g'��������GZE���%���wC&�+E8Y�#v�_EM4�=eG?�,���7�Xr��yK��-�`/U�Lw��T�s��א*UiQ�����%VI:�ea�B��  ��&c�$��ޙ���aF/��^d�ޏ*ֽ��WDeo�X���ǻ��0-��80�f`@5i��&�C��?��4����
8�@m�G�FD����tC��H��J ڽ�9�'��wH\�B<!$Qֽډ�,}ɍm14-��(ĲO8�I`�LS�Bl�<���2��$�o�8�"�듥�yd������jܽ�$�C֍��XF�u ��7�iҺ�O ua�zze.8�a}��V^���$3������HL�m���4��h�9��mBv���4Ȁ�@Q���̌不Ŧ���6��-NVųr�(
F��߆���MH�y��k�E�R��t��`u�k.��o�u?��r�H�B����KA��$(;}��B��l~!+1!��,ظ���\�dՓ�l����TW14���vyPR�u1��cőd���[%�Vyz�!�,og���Vŵx� ���$/�xh�͌6���ڲ."��O�&[��B��L9]�S���	j�~���s��U��547�Y�t ּD��B�``�A
��� �"�\�M���@Fk�l���~@�p��`M�X�U���5���8���1ex��E<�oE���F�i�>&�Һ��H%Cq��pw��U�A��p-���E1B���n�6�p�5��M
cC�3hW�|�����洂)��A$}m���&����G��<'����$�R�}�2b?��	�Z<w�O����P�;�O�v��u!�����V����'�d�k1#'�D�|�GM)�y��i0�z��4���=��<��r��ץC���@�  �j �S�p��¾�Sɠt���d�W���ż��]G�>����(p*J��	�^b�.n���z9����s�<�G{o�����uVx��^��R-���cj�8/�l�]C����ud��v��}���ŝ*�yd�@�Ј���l�t����y"K��^��@�V��R&H\�'{�{9dE�x}G��`�U6�#���1��tC��b�o1����9���}��~���4�-g
4�h��(Wo��l��w��R�7D��z�c��hd�~�[��9�pH� ���g��/w1\8v�..p�R�jd�� ^C0]���g��;D��!�hd�2�܅wl_�Dhri�;�\�o+c��K+5�{���H��S'�d�����L9���0Ⅿ8��J.�(��H��2��B�+x��1�G�z������G�T�beF�\P5�H�@Ht�)&ʆb��=��ݚ"Z���efX^����I/q�kb/�U������<!�s� ��[[ІZ!m(����+����*o��l+v%tw$Q/�F�e�<���-��Q�WK�
��Q���Ct0��'�|cUMu�og�'�vE_5n��Tet*�+?���7�!��to��`zpZ^j �N��+��abیl?�-�}A��_����]8u5�����ƻ���BICƶ�v�a &���v��(N��q��\.�Z�6
��qdY��.f?��3!oQ�����4�zh�����͆�14�_�șR"���4Ї΍_R�@<vļ�%����~��K��b� (j9+0���L����@,��������Xl��i��������ڿ���a�O�ނ9�����B�;lU��w�*V�(D�S��������iB\�NJ�����g�X=��4�G��#�
G~U|���kfrh���j~����FZXv�1��.�|�[�
��q�U�~b��>nN�K
���p�χf���9A�� B�$�Lv�v�;��������Dun|��\ �5h�"�(
�K�&��EzRdt94�L躂��`���G0+�ĵ0�=T��/�4�,e��6��)
��b� +�������q�9�%����=wx�V�V��^��bl�t�M��nS�=8k�mq���G�e+2_KE�G�������yg�~��]��)�BU�R�v�)ƽz>�RWs�=8Qa&S�ַD#�ؾ�����'��\�ûa3;?Ǉ"o"]"��d(���tE�m�� Q{ ��/2��H��8�v�L�b��E�m�^'r�~q��__�`K�X��iT��}Bu|^��2��㙸��d����f�jF��k�x�ީ�s�C��%�X�F�no�p���~)�	��o҅�S�3uI+��@1�?�՟<�q-V�B�|�Ύ����O|�G�@)��f��C�}jZ���np�؄���]��F�N����s꺾+��xCiK(�g�r��д�n�k�`�uap�~���T��r J�`�'���V+/��Ϭ�b�
����U��q��pG��k�T�P䣿��N���'�wǋ�d�R�W���
-�t��(��ƤO�Xqw|��&��y#�
!��Z(���h�&(� TI��M}���E�-W½�\AQ��zR.2|XJ�bh���j$w�dũ�������/)?b,�m��挌�Ղ��M�,���O��팪�:Jr�%��=�օM�R2v�H�=�m�}�ܳe�4{�Ͽ	4p�J��D�rCT]�2z��YŔ��I.�Ԙ��.�'|)Y�F��H\j�"��mj�e��.N�F����Ǽ��N��q��ӒU�׸��g(ra�uʿF�b�ȴ��ٷ>̶5��:���J�Ϲ��ƈ&6�p+���'�ē��Y�
O�hzI�����$xϞxq���J p(�Ź�q�7�{�+��Do��s3{�Sn_����i��	���	4�����h���2z�bi��7S��	�)�i���ѱ�mN
�z�T��".#2Y-w�I�8]�Z3KWn{�z��l;���Et�#��g�f�GQ��64c�[�]�B
�x�H���Q�0yD(G�SV�T��R�he�Q)��U�z�B�}���{`��ڰ�a���Q�`���z�a�ά+]�l�� KK�XB���K�UI�����.�?K	~fMڊ���O5��M+~�\� �#���,��c��'�?�+��Vx�P�v8��A��\;�	�H�ZrGn�&���($%Z����E>VEb�����^ʯQ�o�h-��TԈ9�	�wt��$�b^tY�6;�6�ԅM@�R��/Øtaz;���^��j�m����ҭL����oy����'>�3)�n�l����٧,b�n����#��%���{"��f�l����R�4`�
B��'T+^�5���&��K���&�*G�@PVqC�N��;"�6[�Y��NQB�_�y)iyV�5�Ǝ�Sn�;����j�F��4�Z�E!]ޤ�Q0)یVۿP��^��U��o8V?����OU��k�*�O�p!'(��vS`��>�m@���z�1�������F�;V�3���yV��J��H�1��p�AGm��^���F��b^<�'4��$�0�n�/�j

��1���y9~�Z�n7�,N�pRq�B�nM�Nx�ez~��5LPO��Q���iD]O�6�e��8��Ei4�qmdH>�G�A������b+�
IP��כ�餾�����y�g)���W-=k�߰Փ��n�$�:���n~|eK��i���Ư�l���q�����{�>BB�MFRv�3���� A���qD��]K�U�L����=G:����#����<p�?�Xk��.��Tf�Ȉ�s! �:`S2���"�Ba�o h��/�m�JI�� ��,m�"�pe��.��,�: ����'�=a��)u�G��W�t�`+���|�w�'P�E�l�ߩ�1X�*&UW��Q���Ν������7��qB/D�$o�D6?i/t�շ��G���~mI��5���x�*�z�5r����;C�<&?E��+_���h�n%A��|ԛ����n�U<vHX�V$�9��6�g��k�6�z�#���&�?t2~tRJ�N��v,�a:��Ԁ��k~h}.�Z�
*�*��%���ł�k����j*-0|����9�l:�>�B:�j�Y��m��Y�J9�rF=[����-��ɉK�tX5���Z3�i����O`��]%������kEQoa�{�@����w��p7GJ"�>m�ٲq\�<B��� �T��y�|	N�(=툜_>�[;ܘ%Η�������;���/{���~č�>&	oB?,����i4�/޿
�2u\o���ϲ�φ>w�ݮ�e�)�)�
������|Y�:t��p�T���H��8����S��:��`��r��x�-�)�(>W��4�u��_FR�K���+��r�$E&�M{d4�͸ ��RX�:M��7_�M�.�DճIz.��:�7M`/�HRj����6�geT�A�?9�h��X��x��ѡ�2�}�ڇ�~,T΅͚@��j���ְI��"���ʎ�=[��S���K���Ǐ�B�>�cR�o���II!�P���ߍ���ET-D��UX�BC�ֵl�<��HNfcЗc���=���n�*�&����,�9܎~���Ǹ�A֎6�2 'z�r ���s'9���m6���w�o��ﭘu��V���C9�l�A��]Cq��4�A#k�寜ߥ����fӋ��F���|����qV�X;����T�zM�������W�����]�#��ES�p��ʳ��C�W�V��<�x�mXT�UW������.�4�,��ˬ���\O\�S���D�~3I�:��%�ڔ5�^�L�1����c��)��a)���ׯ�c_�-y��� �%e~��]��|�h���){�������d�f��C}�6k� Rt�J�[=��K���� ���b�X��4ȵ�GA��J(�����/�>���,�2�< �t�1f��=�ko���(5�.�te8���
�/�!^�B�ɥI�I��j���؏z(�:$�[6���p+�|	u~+)D�ӞS\�6��s��;�F1(�ƺ�InNC�,vy���oڟ��t�A$	ֺ��._c�0�3JҴ���~�h��ԙ���$~b�d�O��&;�H>
�|_�wO	Sy�� (��/v9,� 4�o �T��`�*I�gY#�_կ)iJ�& �B�ydO(��[-xjv��_n ���,�:���;��Mo8٢~!�0�ƪs��W<c����Q`)�qjG��z"Ü��k���s�;����yj��g6o,�x�j�yP�_�?�"%�/�������"��
Wh�2`ϊ��"xˑH��N�_��������/�Y!"�]
�H�bd'��sESLH���e��RР7o�x���ȶ�+��
d�ҿ<�&���1C�S�K����1��6���7АE�G��p ~����`���|"x}H�9�� ��7+,��źAB�h���A�{��L4']���r?�g�/l'"g���R7J��{�����W�*&��1���٣�3��;�7S�N�ʯ���5iPg��I�_��x`#��/ۣ����C��Y�fn���.>C��9^���9���:��GF�>p� fV��nq~ˣ�	K�f�z�z�~�P�PT��e|��}�:���̧ ŕ7~�^9N��+�ӥKj��6�E�����N!R�(�I��%pL*�@	
� ���o�BT0V�X(�ެ�̻[vo����x��S�X\���4��=֎��GS�Ԛ���7���/�bS��hQ�4�-���w�~�&�4�je@���p��}'w�>�lm��J�
�'�T��}��I��	-��S�9��_��PfT&�Z-�]���ؿ�