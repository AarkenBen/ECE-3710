XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-�]Rot�&�i}�ɡ��X����&�Ŋt��~Fzu&s kI��L�"�~JV�wq���bw0��%��|��Ţ2uj����Q1<3f��΀��HR	����B.%:��Sp�t0پU�_ NcS��,�BMT4��#�&�h��A^�i��oBc�O�X��=�c��l�?��5���7�Q�g����i�^�ny�b�1
u+9�<��MiO�%9�̱����;]�޴��n��`$ �dP����0g$�� �P�Q���'n��4��?�W�(m��aP=�^<KI�#��DU($������.��U��8Q;_��f�����M)�wǿ��!T�[z�݅�Ub����0e^��\C����=tl����?�#���3�)�1��%C{��[>`Ԯފ��E5��!r%1w Y-m�1\�NWh��y����Sh/���Ҿ�'����꥝���¬�b���g^���b�^!��QpV�;�����QZz=��]�6*#a]���{C�m�k�V��`���_��+��!J�-\�F�0 �8�]k��SӦg�U�'{>��_	]�@
��;��9=�� #q�)i�n��[4^2����{��kz��g�ӻ�&�*ttn�� ��9xoP�F0�����a�oO`�A��l��I0���m�)�+N��ꄯ���+�w�y{*�)�c5�yi��7.��R��I�Dwkjg;�FZ�ea���x�K�)"koaಠ��E�n��Ag�~SŜ��'p�qqr� Ҿ�P$
;4=�XlxVHYEB    1427     840V)���=�d_,#�2��!kT<!���M㢊��1��[+ �¯z�=[:S����v�Sl�ˊ�b��0��20�d2)<��,���tOb�怾))�
f�9��ȼ��V𿽬�9��;��p9I��%$��S:�f*Ā΃��Y6�Ǐ�O�)�D0�ހ�u�^�*S-9ze�m)n�,�M�)�����e����;�;��8@x�9�P�t��IV���A�!Io�]�����cﰳ�)nC*� �u��i܃g43��g��|�q�p�:��rW�?G��o�'�R�]L�懨HK���u�Mm'z��T������>�ڨ?�RLU�OcI@#���-��/���T{�R�,(���|"�y���m��9��g�[�)�_r_�c[����&�|F�ʄȰ-����E����%�|ҕ�� ��.�b�ث �!JvN��)j��<ߴ�K[MJ1�{v� I{[6� �4V^�=[�X�j �َZE��:M*���e
���k ^�Q��?1������C��_�v���U��̻@mMM�a�mZ�.��vX%z9s�{���{vކ �n/=�6�{NtQ2��ʤ��Kr?�ļͪ�ŗ��P{Ԧ�Tjz`��	i�� �FhW)�w�[�p+K꿅�Y�]P�>��8m딃S�Ӕh�i3�Gw֠J�z��@Z�o�dV��g�.Y^�$�)�����9��J����I��ODLĠ��I�s����5C��h�pgmXh	���(���v��7k ٳ�r"�f� ��Vc@�`y�O�\�X����:e�3��������_D9����Pvd1b�p��%g"�1n�ج�W烢k�)]����t�wMP�9��^	"CJ;z����(����?��y�<lS�TB�\�Y��2+�����6���8�����.�R�Y��6pB���:���b��I���7�Y̧��sf�IF�C��6'���b5�R�Lg����
�U��t�¦�$�n���ج"�l�?�!<GĹ�jmZ���:INs�3�%>&�P2ȴ7��,\݀x������#����uޝ���Ȓ{�J�5�8�;C�Skp�*�����'&-!
c��pݫiN�5�`S.3JOw9�|l�G������Dmo	W8���IJ%��n�GAw�ƥ�k��k�X=h������@�=��X�	Z}7��FH�dγ��E*1P<����G�۞����Z�"M�e5)T�Y��=�m���u~�%�DT�8��j7��9�3�U�s"�4O?;@o�pfs�~,ʵRi_;/!�TѶ෴�.�@�ھ����Ѵ����a��`�������?Li�]��������y���V��YJ��i�X�D),��6���M�+��ך���'k���"�#�+��#ğ�g��:��i~��Zs��� �Ǜ�<��`(hW�{��YG̡�g����Ǿa��v|����qB-H,a��B��@ٰ�3��m�E!�׽D�Z�!���k�4Pf���ǀ�e$�7+ʏ,���:a�u=�A�nU�D��$�::�1{w|�` �@��(�s�N?t���)mO~����V<�7�<�<:��ڨA"��S~=�A+�b"��m���X��D�GP���yV����Ld��_� ڭ���r��lS��y+#�r�B���~��Z<�_��R��u�a0����C��[��#�����.鋋��-l�$m��Z��y����.��|{�iL�&�Ef��Њa��|��F��$�/I�`Α�)l�vh%�Wcz��w��䥇0�tN��> .;l�sW��|�u�b�F_��/��S�:��b-c@DHTkM���#�[�
�Bȓ9EC�=�����=��`A�t�
�E���Ϊx��̧o�c�㫀u@�k��(�Y��)i�J��,��,�aq�F����[��RX��sT�SBX`Zh$��i��q��6���`m����ib/������3�ڡ��0Ir�,�5(.cmG_���	R�C��y�A�!'@�Cj������kp%�@�ܧ�
���= 8Q�t������C���X�gi!�?7���C�r��I��/ЪX �h/V�Z