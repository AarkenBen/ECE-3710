XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5�p�2�t��N/���R�h��/%ܤ�9�|T�����hTbq����Gfw�no��3�l�3$7b���*UQ ���)1d�>��VŸ�SU�n�-8���[�YV$�h��8��qNl���#��x�.:�H,<E`����eͤ���6/'M(%�g����qzPHU'q���M�g۹q~Y	�n��X����Wje.w 3?���ցZ�G�z�ȃ�v=��8Z�64R=��/�U����O�VV��^�UyY�b�jT��4��e��&Լ�J��?�����F�(�'Y����׺�a�������Cok�,QQ���74R�Z�MySj��GD�\<����+ �\VTɫ��.W�p�|�k�T�[tr4�8GE�ƀ��F;�����'	�e���@����_��Z�B�N��zBSw'[W}�e��~k������p��[���K-�=��@���76��k�完dD4�n�%o(�Dj䓍V�LzX;��9�GUuV	Im��Lvb�H*���9�J}S�d���U�����Y.�{H����5�[��f�`Б��*��@�d�{	O>�?�+���`�h�[�8��
���C�O#o/H�į��?Ftr|��
�Rˬ����TbD�N5_��Q3��Uhr��.0g���܍.$Y�6c<���^�Ke�?#Bq^\���>��(g�s�ޭS�,(z�hˋ�1��y��Ƙ�_8����1]��#��p�՛֑$�k���X�4`̛XlxVHYEB    29da     af0����m��j���!��[c�~i�?f�'Npi�V9p��C|��3��*�|���>K�%�]ޔ�o���S��a��[b�*Yl�b����e�F�����xHz�{5���&һ��U�:]�����N/4��<�p�C*&����_'	��&-+7�x$hQ�<o��
n^�CoCXӼ��)�����oLm��$u�����A�U�QI�v�����_��&ŗ��ޗ6�҃a=oHkA�J���Xt���qԴcbK	ō:0��;�1���C$��i6^��Ш4�����h�M<���;�(�7a:&�"T _�(���lX��3���ϛ(����(G���Y�f������|�٫0xFÙ�FBg�O4E)&^��c<�c��y�Dq�75��qђ�%p��b7�����H0'`GuV�'�a����ڪD6���Ӿ�k�dB�#2iːz#��+b��[Tt����*S\�a��1<�7F�����Ŷ��t��Z�.,�~g���)�j!A�f�p�����ٲiRLgG����yCb���uX�ZBIr�'"�*qlor��ān���9`�+�dAz����')d}�p������g��v#�ǐd$��o�3����a22�t�=1z��D�t��G�|gS����#:�`4{��+D7S�#P#ep*.Ũk~I���ov&�&o("Uz��/�N�ھ�0���2���<�j������E���c%�:Sf�z��.��_� �X�5��f��wS6._NPՆ�:�D��m	0}��� yy�����-�k%o}�`'3�7�����(�O%'�_�0��_ي>�VR��w���g���QI����ky� I�Ӝz�Ю��Z@�u|\>(�p
,�"^�O�b+����ygJ^���Y#��&5��	�K0��U�{|Y3 �3|<�'�oV_l�~7CW�U���Z���	���m�E<-�ǖ��˿���AT�b��=����rW��Bxc��P�Sd{!CGdL�b[qI�7����v�K��^C/seA�n
���r^c�2;���w�y@<ͅ^�_Ϸ%�P�d>�MN��x�=)�)� ��E~7YQ��P3i"���n^<�i�hY���W���6�
�ܿ���9ҿC�6B���tڢ&*!����W:��6|#0��a��奨��4
��C[6W���֠6�U�q��sg|�똴)S��u��W�A��Dg�*��d"�v�A�h��f!�X�%���o��2���9�I~�ŧ��`�ZQv���g���:9�G������rR�|��LZ�,��7�P;	D[�1�6*I�
��@�Q��h����|M���w�/�Ke�n�t��ɐV��6�YV6J����h�\��R��y�*����{��8��d���g� ��z��E5���O����?�A� �L����S�$C�G]omD3��m�+g�Bur�o;�f1�q����� ��nWA���>�**nR�Рz0�������<�y�E��L܍���h%:���*r�R�-e��I���y�O�*?֣�Z��͜Ev�M����S�R�$�pk���)�_܁��g͵�w��͗ͭ����+�CY?8s��FH��7'���MR����~�Ǳ�x��R�B[L������T����I��]�i�/��������;�����5���D �\,��يP�5�)��A��#pS�,�67"pǥ�b����I�Г�����U�N[f%���۾b/�T�d�0a+y/�v����b���w�=���l�sN�S�e��4��*��i�� 9�q��ҔY��C x�z7!�@���9?ٌh���*G�$��_үbQUQ��E�l*�:�&�����+rx�_t��KFr�zG��\1C�k�ҷ�yΐ̰�=0�ܵ��2�E�`�\�Mp<�װ��#t��=yg��7ڡ{��(2}팿j�.�#e�NM$�ͧ�g��z|�W��Cg��a4N�n��1��E����4Tk�G	��q�|�	1��s���$ύ#�p埦�x��XJҕƜQ�hI�G�m��Jˣ]b�6����K4�әY���{�u$T�M|kG�<� z�0a��~EY�j�����͍�Q�7������V0N6�C�z���߯��ˑ�ȝ�$|M;U4R
�F�w���JZ�A�R�s�P�Zl��m¼�Ad+"�)���2c�qm4W�)��P�*p�9$�uh�G���J��I�S��i\��i��/=�n���?�����;K~]��Ƣ%�`�4#ѧ��>�V�*{~�3�ͯ�
Ͱ�'c� L�֑u1�AAK�h�9����N��B��5��)t;%����D�}�7m���Z?��(3 AA���5,��ErH@�7�3�a�-�:Ɇe@��a�	�KK���">�������W��*4klf~�~Ä`���$؃��ާ�u����Xw�oo�V�������0��|�}f���d�&Н�*��K��g+[x�c)���a>��<Z!ѕ�IS��ǐO�WÆ���a�R��O�Q�8�0�`�i���R��DM��-C;��"�h��eW|{zSH^j��,��\�Ѿ�}8h���L_�h5)��;�ʪy�}509������L����D����QMWw�]�ȐU�g��5}�2Gw�t<��ur��}�+�*&%��5= �@�/���F q�W�/5�#�$Z��! �M�N�U��\���.2oE��Qh�r���y��������f_�@���]�E���e�a}