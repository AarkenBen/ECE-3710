XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l��b|����LQK7|ǂ�����\�{���Ҳ��0�l�;o�^�����Z
�>���D�=�xe� �coF��c��	C�:�ؑMZeWW{�Ϳ�}�ƫ`��5���Z9��9P�mjԿ��N*����0�[b�ə���v6� Z/(z��,(���+��r,��KQE\��$^�D�AQ^e�K/S�	�)�t7��jo:�2�L���3!���%��+\�����8��)5Τ����r�_A>���I���zg ��f[b�#ܝ)��ͲѤ�4ly3<�3W�@9,�����筪ǁ�G��x��27�/�3�g�K���g7ш9釈|��gjW�M�I��d?�Cd�>ѹ@��RUD)�11�Η&���Oy���EE{�?"߾��<��y,3d�ʥI]Ι�"꽊�g�g�
>s��=d�(5��b��X/?xo&��MV[���}�G�
��]ݡ��G�g&>94�m|o��)�oס��JzZ�8�,�u��d=,�k'�w�<�{��8���2�wO����
m�mK�O6�|IG�v��_*mq{���89�1��T�u~��cb��6���������5X�N8W�2В"���j.�<o�9󟤑��ʇ���5*�F{Ϗ=��ڵ�tG3�q��(ݺF��؅NQh�Kh\ε�ȃ�BgK@ؗG��t�εB�h�[vn�uïA�w�[�]��!/ߛ�p5`�uccqֹ�9}N�r]A3��d�|oE"H',���XlxVHYEB    fa00    1fd0m�aK��`��|u�(�j"�7�a�k2o�h;9L������?&3�>x�A�����&�m��'ǲ��,<���o��Ɯ��)�B�U�
�cc5/����k�zCI.�P�cj��`�<hS���j��N��U6��D�[���r�2��.�)��g#��/����P��3�4L�N���� =�$P]�'�g���0��,l��d�.���;z^�֫�ka�����"H�o��#(�(n�ੁx�M��3���Qx��h$�&��1��!>f���ʳ p)n��&�O�܏A����3����{f�oj�4�Hx�B�j{�:�*���\����9�X:�j�$�Ua@�T���tX ��I�۸љ�Bl��7ȍ�@��2��0�i�Ȗ���װWa�;H(�ZV]o�?��7쥞�}	V�Q����N�qeUHn�HrO�_�&.d�L�v��'��z7�7�f�6�9�>�m��;u{������#������@s�
��NA�=N9�s���%m�k@s�v�LZ�2b�}�\>wB	�4��3P���⓳� �eѰ�y������/�:�a3�ɑ<��\�ׂ�϶��P�T3as"�������5&�y��,H�i
�/��b#�����.�GH��\�D\W�ho3��M'M�E,��	���)�vPOe"�QkP��f� �,�\Go�ۊwLU�C��>�:?���?�q��v�X�Q�yD���S�n����v�)�T��}��ȋQϕ��M�y5����:Ǝ�%$( ��.�@�[�[���zf��2�`"�����*�[6f/�Ơ"}al(�X�0��j��*��+7Rd7L�amv ��6d�XL� 7����97�*m��R�[��J࿮7�רz�<��+V �(Y�َݼ ǜ�(���`v�<�$P/�M����SH�N&�X�}�)=��n�!bD���Ɲ��q�t]�)}�5� m>���<F�|�M"�g�=Y�Ӯ�G�h^p��L���[��!�P,o�y��D̉2�ex;Y�=��7ve1�C�Q�ɛC�R20a;��k�M��!��jюPJI�Jw�ىVNrC��{����l�^�������Z�K�G�2����r�C��M!�d	v����_�P��� s!�`�e2qt���GX�����Ϛ6��_��x#Rc�����h�`�i��Sz�H��O�l����z�A�К�{;��ǽ�o+v�������c�S����]��#��I��f�.z�����O�[���^�m��j쟶7=m}-��3�wr�x:�]�:����FV}���m?ޕ�w�.TY�wе��|Z�{b{×�P���L�q�ʃ��+�X��L҇�U�&�G0;;�L�D�\=Z�s��$|�B�ٙ�k�&[�"Fz_"!q��L\Z-d@�����G�{��CS�r��G�L��L����"L���0��9��Iu�`��O�¸x�� �'�ݖ�$я�b��9�հ�+�2
�5
b���	w�ڻD.�-z�=}��2�=���?#�m�Ѭ2�[$�n0�м���ch6F�a�;p�7��M{�uB�}ghkU	\Y�9���r�_��Ip��񡦈�VxS�g��1��!���]�� %����3c !��cj��3ėB�i��_�a��</���l�����@yK㾷�UX/p#���w����ؠ
�_�=6�at����X�p�Z�^��G]��N�"���:_d��$�w�m�a^�QHﰝ�����þp����^���&�,�Z;�56x33:Q�!���c�K/���3m+c��c6$XX�]�a��m\Z#��d����\���yL>��{�Y_��X�	�@i�d��Z�8玚g���b���+���6O��@*�0�.|��5/u��4�Z�t�����mX��������S�)%e�&å��e��h�wT�O�ǿ��
� ��ŜNi*��P:k�BF_�!��Rv�Wa?ǂ�Ņg?c!�L��Dƶpo����?��'4Iۃi�YcE��7_�#Fb�'*�7Me�j���:�{͇ʡ�C��b��bi�w�o�~�λu��Ά[�[|�<hO�q7[ ���Վy�m�����a'��\��E�7ho= 拺��n�u��!g~jW�����$�u8���/�§�E���QE�HF�B 
�(��#q�S���	o�0�#I�QM�I���Z�Ef�m�<2���)�������u��쥈M_�D���	��*!B�O �n4�;��}��3	�l�Bg�e����C���ކ�ď�������q��'�� ���Ii8a)�/wot�V�@x��#�Zq>��qI���\�3_�-��{&����,�2�ا�����Z�όU��K��Y��{]��r����|��H�̶;)TvX��h���5n�y��O��F6+�_'1�q�ke�
�`C�T��K8�
Y<�~�����)�1�fӡ^ė/3L�ڬ
h�{ a��S)����l��.����������u�^h��%�T��W�u*��x���Wh(�c����#k�y�¿�?�z�b%��jӡ�E=�Čf�O�g$����W3���-�HfM	ʜ�'X\�k�e�l�<^�4�x�tT������ᛐ��7օ�5����<F�q�F����������u��(�ݔ�8�.7��%4w���]�h	��|�޽�����Os;�)��G�ԘًXaf�A79��#25G\�3�����8�aǅ�&�A��s�7e<iz���7���3fx�@�T�C��ȴ���>Ҧ@�����Q��tX�	�l3ER���.D�!?<�=*Q7W-���}��1�M�0x�'���۟��8V��B�e���{
!)(ݙ���6��F"m�߷3���dCc���lO�]�o����R׬#eo�)�ĥ� H&�B1wG"�
5$��:{مq�iF���YV>r_��i� ���t^�g�1ļ��	���]ƃ]n�o��B�v��?a���6Ԍק2vP4�����7|��q�PV�;)�6n� <^-�o�Ux\X��ܙ�q	桐À��*~?�h���o僿u�\�ZH�<Ͳ,�t)El쵼:���c�����[�����yX��o4�!y0[���4��f{���9S�:�����Yl���p�[�K�Lz������ko1�so�u�[ס�[�&��Q��{E�'��9Z�����.�R��,�1��!��k�p��f�v�U�����%���C= ��s�_�����˖�̫��s��~H��q�N����-$����	���$�!�^MС-A��)*�k9�:���}��`0�HDI5��j/���P�coC�v|Fh	W�l�B��Y�*qn�=�|����}����*�H�;v,��v� ��&}�ں���g�ԚV�C��(���	��4�ٟ�����F,u,>S v��1�x��4!�7��z�8���i�.�Rg���d�k�\|�r���C�TLYF���Bd�yLR������h���y����k�2X�[eE���D:t��Xy�bv�YՂ��;��U�^Ɏi��a�N�����P�>lDr!��Q�]Qe�0�Q��3���k��ı{�?�]������l�M�e���<� �H��@���/!0�b�m�6cZ��4��C�no�IG������]O���8����m:C ˝�l�2Q�H�:�kO�
�.�W����fiG��_��N	l����p܇��X��,لO?L
���VU�uX�����*��P#(�\����N�f�|J�ȋg/�����ao�A�t��@|�$P"��.��@�~~�T��ʢ�H���w���'�X���e�5*�/�����瞉0,�c]��ƛĶ�f�:���>B
|��-��H.y���{�IP��Z�U�tq��e���O�nNid;�@�����ڥ5C�wbS0;D���Zw�-J����q�]n0�~��e)y����u���.�A&���ݮ9��"��F��,w��־mQ�@� �.7����ϩ�Sg`}Nė�K� �ހe7ȡ�R�;@�7`�H����}�����^Q'��q_m��M�c_o��STf��-��L�=C�]�K)�;���k=����a=ϸP���%)-���І�gX�9�8.M����c'�CutM�</��B���Ͷ8�\��UU�G�� ���F%���<%���,�����h�w�A���̷��m�2
g�ްUL�e�x
>A�E�Ј��yt�)�Z������W�T��Y	��� Fd��+�?:/DQ�1�"�K���ٗh$|�ExiRɌw0���� ٛ������%k��^`8��CN6�SE�h����2��*q�og�gJ�b��X1y���}�Il7&0I�n�7\lRgN��=[_���ϣ�X�>^�at���ro��׃��-q3�c��d�qJvB<�5/�i�Xg�Sֲ/��u|����P���M@	#�2�G1��-��&v��	g�`>a��3��R��ړ4/f�&ݖ�iL��)7>�Ub_����O�aK�]��}��C�Ii!Sl�9}?���4u>�����f#�RR�۠�`i]�`�/~�w���5$���Sǉ[;�B�n�p�yF���B�H�3A^X��k�؅5���3�!���q6I}t��*��cl��|���9��g��2�p|��x4�e�����D��2�О襧z�G�N2ҳ@!R�Z@��j�����ǻ
�myP[(j��R��tO�rw�b}���~d��W}��!;��$����(��	��J�%k�IJ�on�TUU~�XÿD�n�fMT�7�A�z��'�����~Y ��Y��� �\������~H
�M�(�.�ZP2���ߎ���}`Y�'��
	D���m��c�i{�KI/B>4Ϝ!-,���D����`]ٿ+MN�r��gaF�VM�i{�Jº��r����S�V c�Ys�,cJE���QV��td�T߷e�NE*��Ԏ��y���Ѧw%1d�XG�s��u��*!�^�k�E��-ͨPH�Fjc��/����zlѕ�퐜.=63Kp��"��@xM,��i��s,�j��Ȣ{��˖�����/�Ӡ�kXQs`�4z6T���#T,��������4�����e��.����=S�h�R�����yP��*���)>�b��F����޲�Ơ� ���7T*�d�z�,����_���z���
�_ۧ��8rM?�c� ����,��o�c�(�TK=
��p�(X+�-�1�E�(��$���.3��F�e�и����a�q���vs��6���`��)��~ͱ��|���^tC�yl�sR��P�X��dq�ʙ��!I&�=��/��t��\�4�<������t%�(�N��٤���ɶ�ԣ?�m3��Yy���Nt�6�x�b�C�>f�� 7@|Ԕ;��WV�Ҽ"��O>���*�uR������Ϊ��{3V���I� �x�0�Oj54��U�1�!��q��?�0=�j���bNf�D*��}؛����F�I���z�����:��Tœkr���U���M�Y���Y ��5�����~�"W�R/\���U ̊�~�Aw��Z`��<�y�����\�W'v����E ��ȗ�vrƔ1՛��p�uj��-�x�(�n>�_�	hM2��HX�!l-��]���K�b�qX�t����A��^�rzaRA���h��9Uk8��xpY*�\�~�~5+�\��d튈}�D����d��Cv'�bbv (يB�G+Y�G����bt2z�o�6������G���'l�Qe�uv�d*��Ld�:f��mO\��'t5^�h�75%,z4�@���%�w�]���v�5�xk�� �R% ���=����Х�&���E�a��s�e���]��ӣ*z[�jb��n��t��6s�������z}�Ԧ��O�N�ϕ�"��(u���U�a�\��Ȓ�崬�u�4������P�ҏ�`h�G4��_�v�m�)"��b�Oj�)�~�m�)��.��u��6�[4��ӻP��y@��_����\�܁�8}�>�_�rWI��9�[t�%��q���~���p=��O���Ʃ����ⲹ�ç��CB�7��!X.�8W��;�S\:*c�q��F�P�M0��>������ݟ��;��#�B��l�II6qRJ$�+�L�սA�N� ^z0��Ϭ,&%�w���i�Ii�k8�Z9���+��oD^�1��d��ԥ���J��3�x���B�YU|��
��Qj�7N��k���~�\���V�z�Y�,�ʮ����M6���ҋ����?,�+S���O�u�ȕ[B��FM�Cc]�2`(v=��<#&3�X>�/f�`O�~Sxwd���E�Yl��v��JZ��eiC�p��1tnT�v�~;0��3(��B+�/R��]�1�������Iw��2�-��R��� ��Wڅ��q�T}HFz�߯�����>��0�Rd��ƺ*' �V����ū�ᰚ�ȁ?	�0�I�Ͱ�м��w��^k�ao�q�@;O�|���0WA"��|�mZS�a��+�CLwRn��7����H����
;Ԧ� E����;v$�/}f!�/`��g&�2�A�`|	Ѧ�^Rm �ƨ����H�?*�WҲN��v�KZ����vU��!�p%Ԇ<�#(��@��c�^.	Kv�-l���r�ʋ�q=�R!�w_
ے��ԥ�[��g4m�0z��i��h���VCdDD�{t�?м:|$O�TO��iՃ����+��чݾ#�6&��g�NJ��n�u� 5"�2���(J�^�2ܘD�9���Ӎ���cw����!ש.n� G�r;]Iֿ�%���,I�x������O�e�}�{82B=�ق���ԣo���ȿ�����~���Id5�����L�p��ݔ�������\+��Ƶ�K���"�:'�V�!�=� �FB�*�sD�HSh+�Z[Cp�r�?~��4�`�-Q��/�f� ��J-e�����"�l���*B���ϔh���rV��6?�5\�^��u��qȅ�I3�Rx��9�+;��w�]9�� /��r�D��>��1������E���_D�7h�Pǣ�'��A ՗��	�`_S�f�5�?B;�⥠0�ո��jST�	�t4o[���o���ć�.���xѐ�U�oN���O�݌}ʤ��9A�,���=|Q�R@pM����aU��3m�*��5�Z�1��wYCi=N垱G��rO �U�+(���}V���<R��� �wfbqu�&Y$��ی���m�:fC�l�J�yD8��`��|4@<�Q�\_�RKޥ�ۼ٪���d� _�au?o�ʇ��������)Y�[���#D>ޯ���΍�T�G�rl��R�Sc�U����-ה�p����0�b��ȴ"f�u���L���elth.z�C��}��k�6L	Ir���S^pN��1���e��D;FΩ���H5�G:g���;A~�f`�T�$� �~b��o���q�d4�a��N�FH�ym/w��߹�HھTnôAר�g;>s���~� ��Y�a���@��mg%$_��Δ�2��j�F�m����'	8�����t�Ly]�jW�mf��p�a!n�2~��7�:��-�#���'e"��	�w��u=�<��
�Lo���Hwb��ʭ��������T�M�b
����W��j�jЌ�B=�5�2c��x	ǳ�,�%�d�d-�U���z�E��|�����6|��88C7��o��c\��&o>�vr����n�z�yں_�]w|w��CGPD�w{��]���!��-�,�r �6��md�$�Wg!�P[�,i~�f�p���:�{c�����\���Y(`Å�6@�2J+HsB7>=���U����e?m�|o��CؐXlxVHYEB    fa00    1340?�Rbѧz>�AT�3�u75m�1yU�*lɢ��]�ڏ�����"ު�P�\�H��Y������D;k��d�ϪY��+а[h~��&��L3��|O��_jM�0A`�����(9>��^�V�q�xc�b}X���\���X���K;��H��C�ۤo�ll}�<�Z�c���Fԯtn
HW4�{�=���֜�IV��+=��WM
�j��$��O�*�YN}��O�U��QX�I�~8�bH	埨�l�����r�m�'9fy��j|�<\��Ϝ�9��i�v���������fT�b���#W��I�!�0'W�#�������e��D��$7�*�\�N��
��`��3^>�'@�{]iʋ@"��3�h���3U��PG�u�X���_8�}T���R����Db|�t�';6��f������;���44X���o�-��W&��\��[�z�3�m+cl#^�Y��+[�'Cp�����X�V-�+m���d�� S'י�O���'Ua�[]n����
A�����vjG�j�3�B�S�Nr�d/��ɒl���b/�=u����֨��;[A�p9�G}>E{U��y�	�=��Q�>fq�g�=lv�$�����?Ih��C+��:Ӕ��Wv��z"s�]�F����l �Cg�ޅ����K?I��Ϛ	�4=Y�=u��ӌF�ߑ	?�k@k>��I�@x{?J�õ�8�F���:ݿ�h˦�Ӽ��1�p֗.ƔÙ��J~���sBI�I�@}�a��r�D;o�2�a�+!_06��^��߄�N�.s3z��Ȉ=�kQ}�:��_J��N\i�g]M�M Ӵrs��(�H��G�a����t�r��W��P>:���g������#q�t�߷Y!�ǝ�y,g�M��][@<��A^�#�F�7z|@䀪�zρ�(�Y(��Ñl��f�*�T/���s��8Z��P)'�˱�V���
+���nf�\&~i���NӉ�:�'���\�>X�S��gCf*�q]2˙j��48�BS����X����D����>ܴy���I��I}4K�OmH�Kgb�q�Z��@�p$H��M����;M��(���2�d����V�i�y�+�Z�UR�@�,C��7��LY.�R�WU�����}��§�<�̈́��m�@7d��V��Bo^��Cq��6��R�� �����Ùmi9����8�Z�`��n��2�v���u��o��� ��UWM%jm�OL��_�#T�8 s����P5=���p.�b	�����k�g�˶#�]��M���j������ᩭe�3ɩT�l\EΆ+d���0*<�kt��Vs#���:�T���u]^��n��9�=̜���59��V26J�힤Y!�0O�1�2	I��֛ܶH�X�+��P�Y���@�a�v�D#�ς⍩��/�������B�ɖ����1
��������]U��y�d�	h$��#��aj��&��4_�y��ӹ��x�w@\� �!*2�n��f ]  �å焚�Sv����9����3S�6��j�O���rM��Fͪ%mCOa�,�XN��14��e��W�R�]���yh��3��iE؆�~i=�,1p>����T����H;�$u~h�����@����b흠��źg�I�����x�Є��Ǥ� ���>�b�k��Z님 � �@�Iʊ�����,�^�.�,�_Ӫj�r����}9�!3���8�i�����:�kG���H.;\g��9:�8*uԟ+t�E�S}JpHF���vF���]E�=�i�o���seG�������e�*�,��w��$CXn.{U���W�H�_a��fg��� �|��Oā�zݓk��!�;4o�dIُ������y$�k�*3_��e�ZP��qU�Աa�z���Zm捲��4ǋ`B�����doS�N�H̍I�j� �i��2����Qu�o"m˨��⢚�t#����6�_��&h ޣ����E��D�+��Ly9'�1��rXn$����>��NHK6�J����H��,^���kV�e���d���=�O
�aY1Er>��F��E�J�����#O�
�,,� �Q��<��r��L���zb�
ӖDiC��^�v�e��<�Q���j���piQD�F���Ѯ�)���sͰB��_uc�$Zk�����¦�smTVƦ�*�c�#���;=��Ԏ�e�Ğ��5-˔�\���>8�d���+�yC��pI�}�i"�$A�H��c��ԻO��kE�aɏ2r�R&/���<��cB�'ɣ�8�����p�:��ļǀx)Jl2F7��5E�ǒ���h޸h.*�c��4�d<�ޱw/Q9b��yil�q�F$P�ɇo�Z�c�)X��*���027���{����Y���x�(^�uյ�k�M��@L��A�\����l
?ͳ��\��iZ��J4������@�4�;���L����^ǰT� �h��o+�����Jx=y������C�h{�{ħUZ������)#�	�J3p��RA$��-a7b
(8����$�����ôǹ�v}�mV�g.rP&m�M�˲�ȈBR�R��?��J����E�͕ؒ�l��Ū&[.�	����/^�I�I��\@���J��e�"Yx
� �D�
���z%Ga��Ѣ*�s�cl� }iB(�v�b/}�@�]s�ٿ���e��U``-�T��f�8��UG�M����G�,�Z�Z��L'���� �cC�-�~�-���v5˅�_��V0��Дy\0�P��#��6� ����K�隸Es�B�#�,���v'o��i�g��6�#~y��2����Ȉ7�&�+��X-�6:!}!�K��ݺ��,-~��hD��b؝DA�,�_���iU�[���0�-7��B�y�L��2]��[�nwm6�2���M����d�=�ϫ�gw�*S��pgX�
�t�m!L�M�G�����o���J���|�	���M1�PfB|�s���;���R�
�ѤoM,�x�x�QӷF��H�u¼#��MD��V+�[1\�H�f	&T' �����*h��F��>��"�RۜV���,ʵ�S�ʘFg��e�����D�/���Qɚ�����8�3��'�/�igx.n2���_Z�p��=;gM��r׋�'��0-�0I�8�z&T��B͒������]w;:*�;�=
e��Q{_�����+y+T���Kd�+��2�u&"O��=�hT�r�3���X��1�[GY ��[�����d��[�L^�{)s��C(Q��.��'B�Y�Y����',���e��/�a�,�����P��j[�;�$��@�>����8`�`"���/�u����F�a̝5�,uFTF��d�)��I�9��/4���>��7���AU��<)����+"���kW�c���"��o�I��ToJ��q�i����k]E�̔�oK�a"���߻��2G,@�M�Í�S���l��� 1ht����Q��a8�Q���H"�Ȕt��j[P��YZ��ȃ��_���%K�g�k�3��n�َ���	ķ��+��c����E`���Ɂ���'���p�{��41�"u*�@z�g��Y�W}�i�i}���V��HP��qGLoǅȣ��n�����-�W��	 ��e.�^e��H�}j=�/Q[F�v���] P��'���w��F3�3�Q�Y�yƇ�* �b˦����c5��'�2�L�;r�Q���r@$9��B�)��Z��ʑ�-;lI?v������d.��A�CL۝M�J(�,w�E<�.^i�py��00��dD?�w�U��_�#C�n}�];��G����8XA=Z}w��^���Ľ)!�Y6|��CU�6�4��˨���m#�.���e�D�*����	]u�(vP�Wu�w����g�H"83'H���?Cc_�*�Cp����Ӛ�7��8�Y�Id�I��kP����N�����RS�a���6�*V �j2t�+l�a�9,M�t�p}W���?"C�ဠ�G��ݖ�����͞�pjl���"�[P�9���b�0�<�I���úu�M��>�&�6+���V�T�Z**��u�ɗ��X �ư��\2|o�|)*��F�γ�32�1
� �Q�|��i��C=M������X,�}�Ya*��{�Ϙ!����,u�bfV'����/ۚ+޳�nn���$���m�:[�|��3C{�;�#�@���֢���/G!j�j���ˠ���9�9�v���ј'�񺈋��G�������n��Q��m� �;^�x�E�P��<.�
zM���tڟ�X���m�X������0��:]Z�8����+lms�f�ݩ]t��](�| ���PW�� &�6����j)r��e�
6��~��վ"�L�`�B��_���"�pf�Sҧd���~��uΦzMRG2֧�
-#0I3f�6��,A�I���d(tm+��������S�X��$��|ȟ!�-.z�[�j���8xi����G��C�5(Q]6:	��F�Λ:��-���8μ��v�-�/М��n����<���7�pHq/)�;�U���؜�YGkhMvI6��$�L�	sq��$��)wt�Zd�#��f�'�P�����U��s�*+厁�Č]����x�s�iU�$d>�1am�y�%����31��0�� ���)2j��8������gd�����0t.{�4��Ҡ�;B̍wF���r@��R=l_�b!��F�b���c��Ф��W	:j2�&T����+�fʿr�L1�\j�=�@Q���ö0�6�V}m�|(T
I�VUwԗ��$t3%7�飶����O�]XlxVHYEB      e7      a0�Q=�7�s,p�U�V�ޭ���������::�7�O֙��#�]���/�$�@��t�,jKo�+I����hߤ�L�e4�|��c��$�0?pq��O�KP����{:=b�>�w�mGpS�^f�媽x�d���]�~ԛ�G�@�ݸw�D���
�I,