XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`r��	��Uv�gW��=�iW����S�U�9 ��u��C�]��Z8`���A��lH���*��p��s�x	�պ��"FS�У��|�̓�z9§G*y]z�*=UFfJɰx�u
��"����3%5�f��/W:b�y�)H�*��h��œl�v�4�t�O�������S�h�����$�\{�[-�+2�nZ�ZZ�^W���9N��6vx�@��j{W%�}��3֒|�z^��\�oi�eY#2�)����Q�}��)�ߛ�'�a�)Q9�7�����U�p���-�dZ<7ڷ�X`���Ƈ�ւ� I#�?{#��f���&��21��:���%@8�d���W�n�,���6���G�+�4>�0����@Z�. |,U��cU�ı�P.\
�0��X�O|bb��[%��qg��F�M��4j�+��;�i�Xr��˷wo����d�U��щ"� �
�=�e�/��G�3�{�]��&bJv�y�{�s���Zx���b	�kN��҂D)f��v��zO�d�o��&���@{0�|�+*�U�+<��jWI��f���"���W��x${	�SG���줎��e��Y�b��!��,h�aI�t7�B�]��xl��agI��2Έ?�
B��kO#������^�:��j@Am�M�0�YUe1��K�si���4l>˹6���R*"��O|J��W��*�p�|��A��`J�d�����|�(9����9R��]��CA��h��4j�`�J�yXlxVHYEB    fa00    2030{���8m�	���;�ߞR@��Ş�|`�u�����١~���T���|W6?�~���Q�t(�^���ҋ��>b����^��>k����X?�`����Ac�2��R�P��SE��L<Zs�`A��>廬�VƱ��G����4V%��,�Y�̾bY[Q�����.��bB��X���JVڹ�rbpe�\=���n<�rKj�hbZ� �Jf��3\�#K!�?"�8�3�w��,����	ё��Y�����_G�,H�ZF�����ka�b{���bS�Ã������hɊ,=��8mѮ���}�r���@z�V�K+�3 ��:����eh�5�!6�R����|D@��w�	�ܮ������_ޟ�:�U���ڄ��1�O�o�����α�T�	��~X{�홨����ol�ʓoa��<�6B*��ǔ����y~����3�����S��/���@��j�Ʉ������H�!%�����������<F7�93���N o��7D�i&�e@l��F��-��tW�ǟ�/N�����E�)��R��>ʇ?g�����o����~E�ګQf�q�.Xϓ!`�!I�����7�Oc�W��hS����@�.M����+<��kdSAɐ&c�L�{���m �� Y펇sl�4��b��+���^��lg��"�&����j�z����DVq�^b�_,�<�|jnsX����þ1��?�$�G�@י���8y"��"ى���̀g�����t6+c��``�-��K�Z�6 %+��#ڕ��q�Z�$B�����`+�/ŸyOp�ua�P�����_o��� y��|%-�M��)F� ѳž
��t��E��Ucu�ruh|řw��y�Pt	�WT���q�/&�92�߂;@IR5�M�M�J��'��Vg�,UB�ᴣ�#��x�L����~�].���*���SR�ʺ5�>�}Q�q`6©�M�^���p���c�V>�ud�F�A)�%�{�$����M,���}s�ߐ��<�rJ%C5`v��?�T33����KB36N���(��A8��Tǡ�Rh~�2�=�bI[�+wW
G��i	H^��d�hh���+�=���ؾ]���oQY�f��D�����w��ŏ2��O����=����lè�E�x�Gľ��e�&LkY��0e���ˑ��{�6O���0�Pq9��*җc���@�HlvYU{����	�1^��9M�l�ii�S�D�5�Ks���t�v��Tg[\)�ɿ�=�K�m7�=��Lֿ��f5[��E�U�p
���@�h��_��T^6�G�z0�Ef�K,21&��9��+gT��CI����*�����N�2�`�J�����9��ݣ&ؿV#��im+�t�̑Ý
�NgIN��O�1ݣ� �	�MJ�~[-T*&�	���XhD~i�nh��%h�<�� ��~��C31H"U4Y�x+!����>��p`�����N��w$�8H)�4�O7�IkT��^ {�sw,��"��@v������Kp~�>���R /�1�O��s�=��|�S~�����wZ�/�B�[�~�'I��%�tJx���0b-IAg�!B����e�x���u�wv�˵�5O��Z�hFT�>u��V����@��M�~0m�����t�'��\`�B).dE���.cӭƂu�c�0x.�KF��gЫ����Ho���'�Lv^춽>O�g����2��h�6�ſ��m��eTM�{�0�����(O탙Q� �-������{$��#QH(�6��7�>�m�83�K�y���+ԥy�k>��8�2�"�CUEwg����͕Xq�Yl���:c���
ؙ���\���C?3�buQS|���=G��ƪ�����S��\1�@�a��$�����sC&�-T[�B�8}�����¹4�C�#�T!%��=B6��3x	�&, iR�` ��������j�CC��7��A�pq� ��RE���*��4��=��Ğ>����|����.���5C�S�x`C*k�h��7_������Ң@ɜ��Ҍq>�\��U��Y��ɔ�9D�D ���R:���a��|��j�h J!��C吉S�����"��}X����^��9��poL�C�`��
V���Ky�q�r���vI�FOY�v���N_�Q/��H���h5{�@߸✕D]S�ڥ�o�J%YmЯ�;�죒�#�3���m���u*tI���щe5�v��@f��V,��3/}���
%�@�xE����������9Cx����I5X���*܀Ct" �C=�� �QwU��jW sܿVl9����0 �~�?�
Љ�2�����������O�n�Z�r��o�s:�50Z-�R&L���wO�hI��T�o`W��h2�i�a7Ұ+�sB�8�q�K�t���SPǾ��sx� ���#O�*9'̔�i(6�V���Y*�AL�&�Ե�:��5����IWg剮��/�WZ
c�o=Xfr�����-�1���0���9%`�^�xj<�9Y�B���ϦO���63V����g썁L��kLK"eѩ{I�O�T�fk�$Hp�Y�째|�'�h�/�6��,|�+�HFB����ߎ���Lt�m����D[�&��7�)~����b�8�Hrl�	�i�H��,����BZ"�9�Hϲ�gl��b�; �[��nY�8YP�3����_O��,(�opC�w���0hj�uC
�mɭJ��y/ ҆��B�a��=K��)���^O���؉Z�;O�_�
g؉�1h�LLh'���~{I(��S��E`2	Iz��UN	��mu�����|r���f?�YG{�C.�o�����%
����i��������������Kg�,Os�=
k���ύ�Q�,���7kCb��U�rbV�^<����/APԍK��q)�~*U��=!x"D|��P�z�×�*�GM�3^�i�<?N������礶�[�e�o2e�f�˟�Z�Y��o�����O2�Ź�ns`D������C�ANR�Bk����:Eg�u�⒏�㺥��#4@��Y�w��"o>^N�ơ�����$|�=��d�|OiPR��i����$�t�����]�)w�I�#�
�\�&��홝ї����e�ku��u��f4I�J *��*��
�e�u�]!��80)���&K��FW�AI�T�o$�l����-��ye�kO{��4�w��FX(�r���|���iVIh�;2�w,���G������łDH�xis�H��7�7�y����BU���Y {��o�2R5�$O�l[���,x�kK��Ĺ�N��Ȓcw�\��ܘU?+2u^Zp���t��$0�	�;�I��2\f����O�A7�l-{�A|��uq�{�nD�}�<H#�v��z67E��ܲt%�S>/�ؽ �	�_K����#?�C��B��O�.�?�\e��ӽk�4��x����w�ȶ�� ���&�.<A��Ʌm����+�3�uO���ǚ��a�*��0ž|���+���o(����^f��~C�l�U����JǓ Ջ����Z6t�B뜪Ԓ�\�V��[}�	��qy_d=�_������S������O���yh$�6��M�^z�R��9Jz�e�g�gWX��} �#�t��~� V����$G�e��݊���U= ���'��C���ٷz�&��%	���ˁ��/�O��7��cIY��s��;�]���]3J�g>O��v#5�(��zı�",!PQ2#W@���xR��M�_�i�ZG�������=�%��1�"���Q�'j���C*=�T�Ճ���6�)B*��ig��p��u&�2�ws)�Wb`щ|�s��\?Ԝ���X[q���
�v��S��\C��5�ޙ�������������҄* _c
Wn��

>)�#��v�9�m��D$Y1����)"�� �uTV>����F�e���^�ށC:�w@��0�m�H'hT7�-������D�oc�n&�O�&��������n�����.�W��=�<%�Z�a����kg~s2A
��<e�a��O����"�4�h;{�<��P�]�q9ދ|�u@
�I�FXeJ7�)�>=c�:�Q*�x�<����n�e9!��z<��6��R)I��l���2�'�N�Cj�Mƍ�mr�D5j�����{�#n���X~�$��i
��WItɏ<l���C���Gp������m҅��('�Z���5����ꞑĶ�4��G �c��{���X�t ��a�]	3V���4!ۙ���'�b]
ch����b����W�,�^BT3.s�ލ��@�T0�g�l��u��@��'�=ZU%�
�gۘO4����b�&S���֦V�t��g���5w���\�bk��;I�|�Ϟ9�hd��H>�#����T�8;= ��JR���Y���
�ئ߶J?���\#7������j,d��V)C[0�jxg�3�1��l��Z�72hi?��O頠�a��)��!x*mk��F�lf�hE�S�h;GPZR�X�;��M�^@;*ufm�@KH�eR%��哳���5�,��7&��~��-��DۗN��0KF�ޕ�� �G�*���5�Y��(��=ـ�6��� ���Ưd&�L���� j��}��sXՅ����m�����o\��~q�W�p�0�Τ������`����B�U���D�,>ق<:��bޣ���v�Zar�g��KѧrŘ�>��<�|"��J���@��ň�?�f"}���=���_�p����`��ME����=�tnޖ6eĐ������([��X�P\/��<�$���d�U���dQKv���[ J����� ��6q٠:i���T�1�̂���
�bt�1p���"���Ј�P�>��P�t�a����V���(q�p|K	o����%\b��Q��h��������E�[ue��J�l��k]8�U
-��N)�!^��K��A�����aU��D���˂K+��1��Tj��v+�+ч�Z�4���t���R vꇈ	�K-�Sײj�Q_�G-�!�m��$�r���"͇qB��Pc��b���/Hw�޷EPio7�8�<��E駂���#�Z���R`�e����%7`����Xw�+�I��ͺ��op
�H)�v%����x�� twT�/3v��/^�����_��Y%[w�x���E��:�ĳA)�.���d���|{�M�����C�*���HQe;�O1�+̾Z��d�a|���+?���8�yztiE|ù<���ݘ�$��8)"P�k'n���Wn�F�kiAc*�g�js�����dbo�����ɬ��I_�%����\f{�]�3{��?�%�1�Ժ�@�L��j.E������q��w��zv�-��	?����m�Xv�� ��j$��豧�~�������>n�]aÕ��Ȗ�R��#-�>}���\�J�h�:�|���4)��|�k��aT���	<�UdA�[�h,]�(X�5g�[�qk���,9�����z��t��8L�`�8�X�m�Tf��H�f�}�Ѽ����`W_Z��I�-�t��E���j^ފP�'d����C�B�`����{z}�\`���Lt���üb�A'��tG'jw�=B�GZbj��2���?2��B>y�P��K[��l�X+@�f�X���|�w���c��L&0��J�:9�$���GG�g��l���ƹ~�sz+�-샢��I�Z��$��Rj��d�[�����`y�Ð>�:�b���ȗ9����;{�(�X�(�2	����;^��T���n
�A�cC���Q\l� u����')�	�!���<���Ž���p3Ȼ�:�f�KV�LCG�SQ�'�[�!�����J �'H��Ͳ(\�i�V�n��U��4
��)I	��1�t�q��S/�Cn3E��N
$6���y��s�?��^��厶�EMP\Abd_-+�HB��T+J��y��\��Q�`�U�R�ք'7�«^7 Q/��?�	Ei��g�ۿ��=�=R�UE�D�t�m*�bۅݏ��?Fj'-�m�ݩ!U����|���ς@`C,z����tz��7P@Y�->��^b�Dk �8�$P\&����0i�rY��ԋ����¼t��Q�-����C�"��_[E@,OL,���"�u gT�B���ϗ�AA�;�ʈ��ڳtuv�.ɸ��9��U��f�� ��(������{���W�T&�{��+";v��%�����?\:�܉D,#8�����nvOY�Eʄ"�Vá#v.�3�)�QY��c��M���5�z���)��Ґ����	t#s���D�M�u�,KA�B�5���F�#T^��N��^�{莩MP��Sp�/������b�Bk}?�u~���	pÂ�
�1m�!�q+��h,�,�%z��x����d����|�VJ}ȕsx�ݖ���DWy���@��:�=���M>k3�u!�ď�S�6Ρ"h�-������n�褧-O�=�C��N��\1�	��:c���ّ|�J�/��n�qc� �Y��^�5i�x�N��n�Z��jP��5�����3�[R
S�;,D��Us����t->�+�D7NO��������[B�vv�x�B�U��G���h6K��M�QiE7[�%M�H�% �2)E�kYD6y�2!��n�̋�l�^,���y��s�k79Ky�'7V��pdQ@ߙ�������s׷�S\���)�}�.�Y6�V�ዝx�(�߂G	$�x� .6�I�Owx7G��I�����4�f����	��n��ͿI�͈^v}L*����3hj}�v�?�*B�E�K���=��ow�.G�����ا��3�/�$���m�C=7кy}'���b��@�5�o�y�7�d`�zޟ���UO���MO�!�����fW�B1Y�y�������k^"=�,)�Z)C|S�����kX��*&����~
$�6��L�7����}co¥�.~l��y�*^C�����5���;�F��Ɣ����9��3��v=��?["��I��]��?3�*��ЦN����g��bJ@^S�yQ�2?� �^���j�/~����i�X��M���y�����83apcw:$�g;tf�l��"@}��̧���WS�Q�љ+vBOP:�0J�{�������<�-�0 ��GQeCN�74;�`�G�1d��/�2?���愜qp؍�{��L�>&�:�\O�A��8�q螢�=�jk�`k�Cn�0��^��i㋼��`o ��v�YGH�������bn��7G"���,�R�}���Q�"ب�����np ��Q��1�I�X����L���!¥j�<�u�[�Cx�m.�'�,�L��n0 �u����}���e��\�UNO��\����1��Ne�o'�`�������J<�/=���[��c���cr;؇�4oa�����f��
ri{U�U�57�ɏ�Ûp�-�Jc
��5���..c��	�����h�y��x��J� �pXTa%=e*�J1�7T3�:LkBg7����0��w���f�Z�1s�41�X{�'J �X��)��K��\���z�V1d̩�2�Tl�N�A{n�gOy�Oa/�~�㮆jM
�*̐S	D=E	����O��]��=��&���s7[6�a2c�kwϘY�O��LBS=i3��Sx��FĜցA�P�w�>5Р��F��Lk�f�ԡ*�BM�Yɂ���*g��"�Y�@?Ǿ6���Z���kK�I�p��w�aCf�O���n}�H\)H>����@���FЫ��]�U��1��E�K�X\�d�>��<Q_=���5k�!f�֯�������d6�y�(�� 1n�i�ds�4�[��\˷ӆJ�!ܔ�'z��Y���[z烮ϣW��Q�&㎈?�����<�b��?%����7	�:�E�j�sxY�3s|��ӕ��i���92BTlf�:��f�|�-����� ���Of4꧳����,�Q���ۯv�XlxVHYEB    9620     d70���cqgy5�� �To��C��>!�D���_{[N>�E�VSg�z4�I��Ҥ��u0�͚�z�h.^'�N��}V�P��BΡ�ϸ���]P� ګ�-�p��߰�ֿj�k!%�DN=	g�1bvNb�Φ�T�B�hz��9�,��}�՜zs�+"�ymS�ڟ�fn���]S)�=�X�V�I��~9e�\X�v�1���T;�.�uro�#98n�^c�w��R��W����*�֥Q�Q�"i9l�O��=	f�.�����7��:~<��$o������_@�u���R�'�/��Ĝ��W����q��D��f7�R�wmI�Q�u��7G��&t�؟�WK�7�d6+�z	�ֳ�,&AF��)�|7rVwR�{/�5�J#�V�A-<waK��r7:A�CO�n���d��|�98P�}9�~�S ���I�*���r����Im���ܞͦ; 
X&��0�O�ؒ-�(�A�"&����P����X-���`+�+���tVq�P�I��֝��2�D=������q5�Z	B��mJx��y�u�9x48�$�&��m�Ñ�|�i�Ԑ�e#?�e�Ҥ�hl�f����ZlT��T}�����dgQ;�τz��yԇ��HX*��vv��(��W�(
�̳�gEb��㜌mО�ܽj��;֨~�����%�����H��yo�ۑJ�!�{��ɠ��ir�t��Y+%�:g}��I����?�-@]�bct�����e���Y��?}T�����G���-��l��(-�Xy`��v�:4�`oC9 �@	
�e �y�����u��Y4�?Q-�r��8w���ʬFx�?f[�2��wU�Ԧo'7߹���Q�&��������U�	s��,C���9��T�n����t�Lݽ�|�!>�p`���( (������xC��ʓ�Qi�攓\ð{���u��x�c�̓H�|��|�/8��[���n\2�R����޻ަ��B9�'�
���b�m�Nҭ� C��#8b��%�8*fS/q&�D�����|P�gyhb��H�I21j�R�{�4cBB� �'敟zė{�ɶ�а��Af|�i��`�cܨ&����V�R�x�c��⠶���|)�	�:�=���P��+�3�����>��� YM��܌jb�f?��b���׍�7� s�٭?�5�]��������:��K;���d��D�F1���ZP��K<k�Y5��8hY(E�����$���٣��z�v�m�Ґ{^{B���<�Vڤ���[�f�Aauo}#���3T�/�-Ky {�,�&��Y����/,���q:I�exVE���� �4�~��(�N��x�7ʭ�j+���	�̩ �'$9��GC9�ҽ�3�q6��
K}N�����.n��LރK4�}O��}z��`
�N��c�����+4�55 s��ɇ[�WsV
�g|@c��S}��ؿ���Ko�r���JTʋ��O��8~]Xm��}�&7�=��C::,~ݶ�-�m����iB�V��8 �w�&T׷l�#�j9�GfA���P��e��Vf91=$=��ܻ�rlԦ�{x��"��ek�2��(6�g���qq���I�Q��3��9���%��g�}Pj���G����ly�d��}w�H�dW-��UHD$�o[��e�7���7�d
���`� л+�9����fD���؏�LV����iD]�-��n�Q���w������v.�����tI�����%o�}X�~b��9��|�t>s��>�+9/�g���Pd (�5��$�}�9��z�HC6ROM�j+	q�!ݙ`sR�Бu��^>H��V�۔���Z~J�!�7�+��>J�8�	���,��4�Iv~�I�8��m/�k���?����~�$�S,ho�\K>���RT"���o ��؜��F=�M[�mM
69��&�����{zt�x�T������{�<��N)�
�O���뎙�������1��	�X�~�z�D�}A8�1��u
�A*��d�!�Z#_�UIMqo��>N�l�%Bg�,�4}{PH��A�����1�W�udfm�^4�S;dd�?��W�A�mm���	ϵ܋��{�G�=�Ea��ŰT��ܮ�;����p��-â\���]ʿ?*��gw�<�&H�Ջ_ ɩ��<����Ӡ�䥵6w�>dH��ڛ\�mİ'&�����+.�@Yjō�#j�q	k�M�.~J1�Ç8��6� @����#�Q����/�d�0-���.�E4qI�Ks�����*d�;!W�jfߝ�~Z{�L`'��gvo�*C1|�H��l|8����R\����?K����<�Rv����� l0���zf��{D��h>����D{��O�h^A�%o�9CӸP���S�٦A��taH���[��,�O�m	��5�� z4��y;���|R}M^E
y���Ṃ�ܽ�T��Q��ǉ�X�V=��.�@�Xp��`L�f�`f'�WDݽ��J�u@�7��O���7K���8i<�,��twh�2����x�PɴLp�>�8����Jz�3��x���Ϩ¢1*1��P��-l�"������j29#y���G���&6Π1]?�����f�@V ��H1t�n�x4���G�AbH��'�7��T�Ȉ$/#?!in�%Y�*c����/`y�9) ����h;Rsv����դ�ዶob�'Ü���ρ���Cџ���Z"�
*�e��4��¦��w���� 5d��m����G�Za�p�~, D3�ӝ7>��=���w@�����W4��D8&}���Q�lq�iJ�Ťڠ����ر���8���Ǥ�[�(C�@��(�H���J£J#E�
�,��a�� (�Wq�Q�e4R� U���2��@��jv��K濕r�%pǭ�j�צ�]��^���\���-}ܝ�x�s_v��˥à��'��vW�m2p>yǊ��h�笛pA"i}�/_�����;����ZO��O[Orɼ�2b��^JFL�NG'�\��ñܦ�ҩ6�i���۸p��e|��4WBl����(+���o��}�K�n������-LCA���b��I:�*NI�?,�R�r1C��_�P��F���Uҍ�,�*�R��Arv�4% �4��*�B���4������>P����F��s(�|�����L���A�B��N�X'(s��w&����g��l�H�^BۻP�>�~�wl���Ȕ�ƛ0LL{����D<�I��}�T�"%�W�nuS(ΌAzoh���ҶP�V���A���zb�^�Q�߀S<Ɨ���<���ۓ�LN*c���]�ȣ
��
V�R瓧Է�d�w,0�e��SM7