XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m����8�߱g���J�����8i�wg��(�@�O�V��iZ� }���5`�IG�m��j�k�`q,y�K� �푰��Nt-�GG~�f/{�)m.��񩘛���y��~y�K'r��1&�"a_fn` ��V��C�9��бq��q+��1��/'3���t���W��3ix�H /;-��l���h|�ނ8Vq�'O?�+�w���tw�+��BSCs�|lY�e,:̾�|/�3��5��~K�R���VH���5dOf��'ϥ�q��cΟs�~?�z���-ߩtaM�\��(�� \�88�h�3��0İ�(T����Aڎ`�G6���יH���י4�𦓸R���z铴B��I��ó�q���Qȧ�3]3�d�H���rQ2Xq5�)"����}��q`��:M���ֲ~;��8?hң�B]U�T��EG��p�M�fו�nJö2�|��N!t�$H�	�f�Wzk�R�A�HF%g�Ϛc��d�l �Y�7���ܸ���^�����7�D�M	���긐v�$�d���ca��w���6���̏��m6��%�7�����/K����-�ir@�X���݈&�7���A�m�b��Ii �ݥ�Z�4Bԕ1{5N��zrD"+�
�$����b��)T�#�N%+��Q����2y��E��.�Y�v6��R��Bb���L�k�Eァ���Pb
����h�}ƣ�!��jC���%�V�Uí��cv �؁�`
�%���!�Qf]�KΒ[XlxVHYEB    fa00    1f80dǩ�<3Z�����\:��1|k��x���4D�r ����������ޜ+~i#�ݪ�$W�{���?��nWa�vz�RUQm(m�Cq�����1���,�sg��A%��D#�LnS�m�@�L�k�3�L �4�9��ę��d��]�(g�������A,����	�C��=����%�9�`��y�W�wLs���;��אZ�\Y�M� ����	$�4X/�H�.�~�s�Ӹ�TfL3���� �.��x�O�Rꬡ�x�1����A*��M+'9*z7��.S��	T�-��+2/�F%�@?�􇺍�U�4� ge|��J�*�v1�@�{n~+�~9)�S�<[�V�SRC!>Ŋ�������eir`��B4���4k>�ir�<G=>��T�zj���ҿPD�䭊Ʈk���5ƀ�)���D1%�!T|4��NڦV�~�O��!}��SI�&��ՁM���&B��d��`��^�ڿR_k��㸅~��]�oLK(��ĮJ��S͋t���6��Ǵ�$O{�ܦ�X�zB��*�ѽ�}:h�C�T�j/T�����-2e�|�%&�D-
rw�������J�A�F�,2�͐��cz�j1�[���l*�����"��y�#�-���1�|�ҁ��keu��������m�;��F�:�{�4��Y!:�oc����� E��z紩����
��V��*��e ���/$x*�IΎ4��`�&�k���J��,��Q��-K�
@�5�Մ��n"-�KQ$c&/ƪLgJz)�~��-W&�Q�ǃ?B���h,*�~Y�$�PV���.�]\�:��)�l$�����#o�e�k��K0���$e4u��M�������2�JQ>>�mL��m���΅G
�#J���1�g�p]����S�(���r��Ȳ���H�� zO�Z�v'F`���=�I?Y>�5#����Azdda��Z�в�~i�����@"�p:��.��Q�J2�zG��~�*�j
`Ώ����@�ݍ�G&\W�YP�M���o��s��X��/�'Hr���R�96�����(
"8�ve6�Q�HߡU��k�aQ�*P��i.죚�%Dc=��a��/G�A�7�C�n����s?�G-��}pr]'���,�tŝ��_��2j�Om��e{C��yc�æ��/��Ĝ���>���[t�t��xָC��v�٢)_%|��j����Zs�Q�-tAN��T��O%��������C5�����c ��=U;%똓zpM��9�G��4
�_A,r|�%½뢓�)�A����9Wm�J"�e+,��2f��	�P\]����	T۳��	.�JEF�	��+�����|)L@L/�N��2����`)�q�n/<P���S�s��������'��|u'h}�=���d�l�O���g�o���xʓ�A����b4�]��&�U�ΙLҩ#0�s������k�OlΥÀ��<�y���ji���r|<��W��d��
������=�Ш�3���?���=��T���Љz^�?:�I��\�C�N-�e�f�9lK��a9���"��ZΨ�����Wۿ4��Gq-�3�{?���8h�x^���?^���}j�{��G�����GCl�{��4��)+��>¬(� ��X�z<�3Y"wy�R�a��4w����͍u4-R򲪈I�����iҪv��< j(�ys̶���H�T�8�8]�H1��kKY���:~dw�?T,��ܘ��i}�By'XĂIFW�ԹL6jx��۵W���T ����@�T]�/��,��/�G�������5�/�y�ظ7�~{�BOI��p2�a��	�v�w��sHj)8*E,B~�|�3�UE6�t��a����ጣE�0B4�"Ϯ��^�Q�bR4o�'M{�����7��J[ �MF��B��\8�)�h��g6�܏|��8�:���DϞ�d�ڳq���=ei�杔���24thH�:D?�L����ᖖ�v�/k��\��9�����!��DL�"���t��6=��s�;!Ĳ�@K\�Ϭ?���8�A6�ӡ�N�?��D�eS0|)�9,6��*IS��?�����㦰<T��zb%��_���P'>+X�{��)�E�.�/�^�ڎ4v�%6n�Qe�,��S�<a���W}:2�8�����vL�gi�a/sxiލ� ��!�V�_����P�Lo.���2r�uR�]��Xe&�c�[�M�8CH�Π�֋�9Z����c�y��ah�dcPv�Y������w�]��MK���9�^�K!]���0g�=N���$�Q �� �(_�u]��M`!�jF�ur�>J:R"�(�C>R�I�� �6z���g�Vy�=)&�[��%��㉅=��K3HN�(����J�V�6�r��e��G�ڍ?\�a�g��T�fu��@oX̶9��y�DQI����@T�ۙ�]_����(i��J������T���uh�0��Я�,��W��-��S��
�|HXAR�����j~F4�3m\"洋�&��L�T+�?�ګ��\�AF%�C����En5}��c�|�\�Db�b�ݼU��~�7�k^� ��������>Z��R_����i�#N��蠔�hU{Z�y�"����;���U����uԵPx��R�m ����C�a�iD�z�)�2b�:,�"�Ԁ��x��}2F�Ʉ=����U_G�A�p ;q�2�E�H\�NܑpV����ʌk7�f�*�_U�֗�>���=$J���ц�6�����pV�����?JN/�\�����Zs_�&�b�cy�[o�鳮�4�q�c�ڴS��d~�9����=��g�i�1���6��&�Q��?��.���U�kS�;��؍�R����_�L����(��
|l��Gr9�/��:u�U��Ɋ?=¥�ܲ�>��Y�29,2�!="c,KSm���[8����.��	���Xk�,�jC����x���N
���(�q�U,ξ�S?&�]��a����4X5W���v��Ұ��+�i؏���0�F�?>,���)�6j���h��;��e�hMvL�
��m��^s>+2�~o��y*@5�4>Iے����r�D�l�E<i�K�C���|�Ҫ9lXg��Ͳ��mC��;]t>i��ܸ6�?:'��k���n}��A�/�P�^Ɇ��[��]��<>�cw����PD	d?�D�x�g����H笕����Ǘ���	uG�O������\��@����ul��m�1�1c�.�Qre玔Lj�V.B7�ܐ5!�*����.��7�1�~��wJB�<ܯ"���W��7X_�1��}���>�I^h���T�aj�Wң��FE��;W��]��Ro;����<�/T�<^!
�t�&�	k��k��|L)Gn�h&ʍi�c�:�f�%4W������r�%�Xu�l�>jLLy�W����$`l:T�sU �oS�g�m0NG���_ Vah�J��9 2|�7�آ�'��]��>@�}n��&��>�o��.�4?P��Kt�	$+�]+v׎�f�ⷓ�6$\�z���/��y�.@�޽̷<�����1<�k�.6��qa6|�$���D�i���Xa�y�aT�͵��"�2p;]n��X������UoW���O���])K���)ʺФ��IBY{�r]��А	LAf��W��G��,�e"�D��ׁw�T7�8����f�����7M#�,Z&Xx���� �$�J�����Ī�~�2jA1S� ���&�2�TT����@�qf/��c�R���<%t
*F1�9���k9��>z�m��'$���5cS��o�Q/A@�k�= ��U&%��3
#��-������h��π>��+|���H�)�f���Q��B
B�/�w�+���`��jx�#I�Tŗ�j�R6q|�^�3rz�~}sܞeEG����c!���������!��[�2�J~�>���C�&���=�2l�D�DB��kI�^����1�^�Z?��[�jd�I�\z���=:J,]�����kGmxb���b���G��6�C_�B0�f���˧�ZY�?�C@U=�yJ�l��
n>ȇJ��pǣ)�pS�+.���y�~ [�r��8i?�P���s�1�U�QQ��g��y��OD�XO��Hߢ훏��5R�	P����{���ƒ�s�"�u�r��yYO0z;���o
R������e��m40����ZG��<(Br���r���>X��p�D�ON����h����g�d�~�Mմ�a�@�r�?�����$K�=��ʓ ��i���/�)����l嚸�n1Jv�˚E��I�C(�5���@t .ό5u����xdа�>�07<[dm�G�a�?3cw�ZX�]�;�v�Z[]o����P��Z�]�(��k���R�o�?��4>��f�䝻��%��|������h���u�M�ոM��X��dȒ8:'���e`��]�=���Mѓ2��|��icP(��^FV@��e[xg"\�뒔9������:b�mI�^�����
�#8�n5`�>j��7����P��p��0c�~~U�|,f#���b����T"	.;��<%��;ԡ�$��<��R�̸���$�;�s�!��7���4 ��Ц�"y*Jb�W�aXl�bD
'�[+�4�T|L�Ȏ8�V9b¹hD#L�Q�
��-W��	��'C�-���|���7ݍ�	����|�&x�J�V��i�݀O����ȗ��U�I�C������F0��m�|��H�Z����܊�%�*>�6��7Y|��Suw���w�2A]M�X��c��Db�[�&�j�w#���I����]��P�C9R��.�����kl��+���؜H|stb����D�d-IQ8�������8�oMY�Z͘+�JE)�'8� 	ǝ� �C�s�!�d��@s-U\�,�V2�vb�t���Cf>B)v����PS�Nf��V:OI>�5��j�Z)S�K(�"�?=�+q�X$���ɯHٲ��{����?X�j2q!g�A\ǉ�:Kܡ�f��"��f��n?��w�f�w�������Y��?�wE蟋(�u��oj��@+���Zk��|�4�	�q5�t X6jd�э�N}MG�.�WHj��!��ɛ�q#~�y}N��M���`�q�����CEw�_h'���\;����Gp�r��F{,%�$ws3|��9MK��P�q?6$�J�+�90S˺���޸$�T0R(R��u៦��\�Ƚ��a�9E$�JH_���
���y5�P+n��e~����Y0�]9!ǽ�gǂ�p��V�w%9�u��1L�1ɝ����?+@�G���oM�tX>,0��¦��"UJ:��@dp]���gu>��^4��,b�O�t櫽^W�A�7>\�ԍ���	��%���9Z���:*:�����	������LU�O�g�ꌓ�o��zk�E���%���}��0��}X.u
�E�Mv��Xfd$W$�%;U��{0������Y�����6�=8���Ԭ$i�w �o.�"&`��A��I.г�n���}�q��;]����g0�K{K��������� G���Y�|Q	"�m��#qبiM�tnn�{~��N�ڷ��5�j��*$�6�����Rt?���ϝ�:�]�v��M��9����� =>bBv�'�nW]���A�[���'��e�g��i���~��	zT�@��ȯb�Wr�c�fBw��e	�{ꭡ|3�J�:�	�3j3�Mc���D�I�s�L+L�m�'{z'��Lo�j�~��ىm
!��RHQ*�a�j �7�ccX��\o�ܵM*��k �-5w�g�l�s����������(��ht�F��J[겛��2�W�ƿ���Ëf(Zy��@Vd���M����ϫ��\V�r�kȥ��dܒt�*6N��=���m�x϶�n�QDlQf�C'�w�;��us?�*��b�}�+��Q��)CA�X<A����U�ɢ�ڢ�1vHu��A0����B����:H9��lP��$+Ӕ�>���B��	rѓZ�ϓ��B7�4�ޣD�}���W�-��F�]hGm&Ū��g��.u�L�6��<Ύ��c��s�Z�
�b,��m��33�5T��q�b����&����2�M'�֖Ĉ�y��]4�B'��J���,d��p,K��nT�_���x�:�Nŕ8C�D�=I�]9�`�	��Ώ�
j�&R�$�2�b
a�cVIj?E���z�ɣ
K����o�K�x̑��9/�>#<v:�{�h?.YUM��2��vWsC�X�X�Dr�)n����?a��-Iu�'R���˞v��kܴT��4&�Ҭ�8hژ�Q픃EC��7n�a ���tjt�3��7t$��C�����[�Mf���!�-	��i*p��}�����ij�P�ݱ!Y<��!!.�U�Uwv]��v�)�E[��.)�I苙���󥁗���v��m%����EG���a������m�Έ5P(kLk0�,����I�Ȅt!�U��L�.�~��a�"">��7����MS�-�s~��̀��+�2�Qa�,���f�I���y��\p��:�%��ji��fc���i����Ͳ }�b@�D�o��ɶ������]����=FW�����l�6�_zr"$�<������.����UG���Yz׋l�8�$�M��{�>F�2��=� sj/�d!�&��t"a=�8�7�_{8Yb8 Џ���]n�x��uS���0�+����aA���Y��wLʳ��4�鹖�E�n^5!��>~�{K]�
�m$t��X��Pd����H��^���8�85���0@����H����qO�i�:<���w#/�,�ʎ��<tfP��#U����dv�Cf�M���!�l�ģv���fS7�0�S�G	��&��gE)�ƸEOc3#���6|��pRT������_�����,B׹�^�%�yN>nW��|u���Ym�6�-���cU�}�ˆG��{����於f-�M3�+r����f}μ�`�;�&�`G
�Z�-.5>ȷ�$,�6O�W�67p�C���ں����N������KfI/
��֓��s}}���u|5;lQ�.x�q)2W7��%�ӊ��V)�|M� [o��'	�H���>�>�׺����;�QICg�
eCb����{t!�[l��"U�^�~87����`BI'�W(��%) �_�� È�QZZ�N��,B����͌� ���ZFK�k
��s����BɡJ��y���e@s[�!��wI�3�����۵R��S�6"L��"�b)H)�n�s�q�͊����J�^�8�Fh >TWa]RI�3�N*V���2�|�आ&B�8,ٟ9s5�������Y�v�?O'W����qJ�'�1:+�N���#qArJ <�A��ٽp��{Ԇ֌�Ya�D�ʁ��⁮�X�������u*��Z�4G�Ӆ���.`�X��l"�� $o\�,O���L@�����<�W��p�\�9MV���pg��p�h�!Q����:
�s�>�D'E����`_~��4�v��S�ښ����Ϲ���!|@�	ә�ǿHT��g���f�^�s����N�%ں��=Jȓ�S�p�fN�Kl�3���>�a�s�[�.,�p�kRK�rjR��m#UYwY��|�6��B���ȮM	�g���$Y:c,b�xHe�ϋ}��E�D�GT<�ijUDT�d�J��\}�}����bE������X�)i��Q�v=�W|L��ک��w�9����)��ܑZ��L��Wm���VzH�CR[@R���������^ �<�\�O�n�G���MŀI\��%P���m�w�����~J�n<�_du���S��i2޲�tk!��L7�A�w�}XlxVHYEB    fa00    10c0G�L�إ&�ɸ\
�Q��lF�y5L��V!Y<�o����|�6��\<U0���q�Z��L����lBhEuN��>־����PO��IH�F5�U��Ęt���xT�8@{>�01�e�v �Bg����?=��� ���L���.�ҰD�f������Y��WKu�\�!��yVYu��]U��ZM�4��!C7� 6��_W���]�qX��r�I�=t\#�-�O�tt���̼�7�?W(\?�'�Yh�,�)�U�۴y��3�ƼP�,"W�"����:'�w���n���;�	�l�^���i}����,�T�y�QrwY
Lf���A�[,Ď�0�0sG��H�j*o�QY")`�������bڜbKs�(g��=Lփ؍�mm��8蛌k�*p��.M�9;~��3����O��J�0�x����z:@��=�҄ST�ϓ٬�r���gW�S`#x�&Ѷ��k���ʢ�eKA��ri�!���~�Y�J�$P�)-f�~1���{U�A����mc��o�z��o@�ޑ� ��w;�c�쮛fǤ$�'+�����VH� �E?��97�mt����S��[�}�3�;�M?y��=w�3#�yg�c���=��񅺾h��vX�=��&����n #���.��@��7�m�;�(�jZá{g �$�����s+���*�罍nVFM�����	�w����r�p��=BZ��i�~���.���J)�4f��"\�vW���(��a�6��V�0�ԓ�O�h��Z�
Ny,˥&C�������g�];/*�;���$Qϖ���R�Dà�m�8,DQ�[�/�cs�\����q��I����4��':���b}s��'$ B�G�'���gN��D��ن�a���pq���zz4�<�'~�f@;,5"���f0)���ڛ�W�XS+�É��g/���g��H��Ds�_Ҥ�We����(3Ts;�.0���Nǁ�I�WYAO���y��s��b�5�o�k	c*R{}V4i&�~!��X鬕����Sɇ�a���L�Г24�t'*�O��!B}���\7���k�4������!��'�)���߰"�]/��y��"F"3���㲱�7ƒ=MKu'�`��QMϛNY��;���K��.e?��I�t�?��2�@ؙ�S�1����O�7�tS�D
i�l�<��_F�YIÂHÒ�
�.�%@c�����n.I�)�b!���N��\_0�5U������ߑנ|�"Y��֌��şs[���H��xW��+u���x�*?�[Q�p�v�$�A*�ϺY^N����t�M����o��s�E�^C\|�W�Hb8�TP��%_sӄ'9��gS��	�w*�8�3s}V�Gkpj`2��/:�Hd��fz���^��I�<�]n�CQ�Wb�z��( Ұ��6�zӏz�Yଗp��v�Jq���@�ͩ���&ʘgw-����r@���b�%�e��_B}cw��
�y���w\1�Y��p����6�5�,�v�c����.��fE8� �i�f�KC#��~_�����m��x�АV�tC@#F|���m�ىRg7��	��3�r�L�"��2��Zh��ꕁ�K��>3��F�x7�'�ک��L�U�r��P�����,O&΅��Kمs*��N�+h���������R��'��fW�8-��P�/uΖ��d����2�XL��D�Mx�[7���$�3An	#F�ih��d��ppv����O��+r���F�[���N��J�R2����Z{=i��D�8�BD�+�;$f���s/
��+zuJ�A�����c�n�mO&��=A#���lOl�Đ�����NR�Q��a����v��\�A�c��E�G�4!I�x4-{����\��`��a� *o�歆�P�иT���	�7K�v{��@8��p�@δ��c�o7�����D�M�8��(�;���wF�꾛�at˔N:1�hp��uS��ʢB{�iN�<P4yGS�f�U���B�Kq�;�=<������<ߚ_�4&��5H�Z=��vHv�[��WK@X�Sx�:����V|��"���v 2�I�3�G���A��7)*.�K�a�RrA�4��
�^�JV��@��\�Q>����5Db�jJd��tf��Ή��B"}��Nv�7ͣ �?�s=�^w����j���p��}9c���7/�֊x�����s]��Ո6UO �)���A1�u/�'�F#c�x�n�8���%T"��f
	��%�6�A��ʃ���c��cl��և-)L��pS����3i�� �0���Ѫ�4Jڤ+(���9v���{,X�%(��]�Jd�f�OA�m
�,	��P�)Ӫ�@��|�'Üf�v'ICf:�9�*�;[�$�uX�� �e�����W���$��]P��g
l7��ɯ�&#����m��fz%�>+톐q���,*鋪����������1~��=�� i��"�ܣ�i�D�]����~� �]3L�U���6����b�n/�ٻ�Bi�GZ)�R"zw{@�4��Q��E��/�jPl�օl�I_�	���1*��Zp�ʢ���;:��z��̘;[CD:O�(�=��mb�C�R��+$(Ɍ�"�m�c�W��X�Vu�5\<�����~?�uL������Zǘ�x�֕��u>x���f�/�N����Fw��{�i�`'\rK��q\*	bY aT�\���ť؞��2�����F�}-��B����c)��u�J����);����M�>y�62U�ƄM�@�'��wBL�Mny3��M�-���;���0�g�u���ܹ��?�U�h���C4���JF@Ye#a0��9Y	�.CJ ���J[�'OxH��:�6Dyf?^��MJ��dG���&^���ǰs�(����d��-��JH��c@���mb���v��X+�E+Nj��ĺ�g��A��M��o��Ĥs�nߋ兲���7������D%�j~L��ۇ���ҳ�8m������}�����^f��<ܷ�e]��%%��X+�Ӵ����A#��VJn���m��g��Ѣ��G��D�H�
��X?�y��(��&ĺ�S�+J_U��-#�������n�{�MS�1����ᮂ��|rK��l��C�����P�R:a����Z.	}���B���6tE{.4�f�<�FzS5���A����1oJ�=o���1���zY���ѨgN*���W	s�X�9�}8붰�n��<�Y��4��l$S0�A[msE��K�^op�=�b ,j
�����zHYX��ePy]���?�X���wh��ܻz�O��!1�r�b���ܯ2����o@w!ٶϴO1d7z<���Y["ptx�C~�#��p�+F�-��VCT�����a�.63��v�<����J:�.�_�[�� P�>�_}��6�Y=]�ϐ6Ek[٢�y�uAy��$-��-9���5nf�Y`�-��L%�%1�<��DC�]UO�M-b�Q�tN~���CFh�&��_�p��LR�:o�x��}o��g���[�Y����Iv]�CF���I���#����/0��?b�9��'�}'8P7I`4"���Y������Os�x���d4������8�9=l=�A\�Ք��8��r����H0�4�� p�)��Wf8ӰCG�Ʉj޻cji26H"���;'	�U�?	��f�D&^&�k�
�u6f~I,������8Qi�b�t!�0�Ai	�;*��M��}	-�o�c�i�%���D�ci��@�P���괵-��w���&''ANG�M�L�(d6,Y�F���A���G��!j�͘��q�Te�h�V�Y���DU+���\1��΂ǔ�����F�H���<�5a��C�1��3�b|�pW�``_j�$6h���وl�m�DCC�2���Q��t�	�&>���!܊������/hj�L6�����Ii��:�c��o��F���3k�PE�%�|��Q �xtn��s@l��D�^���jMC�w��~6��U[T��1�P��[Het��5Aq??<S���<��%�>V">�3���ͨ��=�kY���� ue�m����׺��I����,͙����7�+��L�|�I�o��k-x���s���ɉ��"���`\��[Z�mt���I���6�R�?�z��'d�8XlxVHYEB    fa00    1140�Z�C�	E/7\�������s��H�����;��e{l�&jn�T%����;0��6mU� �r&P@�D�h�[��
Z�Jܻ܅R<�0q���m�8��Ic��.��?���͙!�0N�ɥ0�rJ$�xXX�=&rSW cL�� ��@r�}2p��[=bCZ�������/=I�-��4匂�����(Cl?3.Sm�z���{�O/���3�|�N�a�K|��  �Ff��8�<}X�,���d̓���$���
�8 l�-�o��-�[����t��F�f؂����҅*n5��:r���D�O{x=�-aܬ��mp�v35�t���
>N��3O�6���D���LO'���C�G�i/��ebANd	�����A��jPK� �PL��0.�]f��i��Y?,�]I�$nR���ߟ���=3$ŷ;���,f��/�ex�<&��X������[���4.��FW�ʹ��z�3�ԡn+E00�,��
�5�z%�=_�`M4��6�u&��C �21F�b�\�FK�Ԍ��6�5��!�uC�y/����?5*�������p�t��A�ɖ!o��t�
��؂t7���!�Z&�
��N��t^z��w��g)�/��N�<�j�p6y�H;�On?]�Պϗ�YࠬlVݾ��㺙S�մ`�OĐ=gf�ͽ���[&[��q��ԝ�"hb�������m��Ag��,�K�/�c�H���� 'XF^̪�(Yǆ&n�=	�D�^3z��)3O�b�&��ܡV���>9	��c��,G��	�6�I�5vt�ӱ�髧�`�G1��Q����74:��ԑ�Oh�GR�8e/�v�In�>4�Bu�$<���e�W�4�=�3=���G�����f�Rw����S���0���\�P��"2�l���|݅
�x�I�Ru�CA�d׷Bi �&Y��Ǿo���<PXUI�tz�q��\�G%�~�d������&#C��j��g�q��^[�7��B��"׍U¹�b�/����cת.e�z5�)�G�~��Ā����&��F���1�HQ�S:�"�+��<���"���yeU4�ȁ�X[���sl��pW�x,$ �E���Oo����.3$�M`F�"#�[��L���o5���d@ �M�h#��#D��̵݆����^1�I���{}V�5���LcG����f��	xG 4F>3��B븈T���x ���N8�7�f_��$ɘ�])X�`؂~!������<}�=tx^QtI���q��MI��"9��&j�h�R���Ռ�+wxu[��Z��U��.� �����;���7Y��W.OȀdO	zl�F�Or�v��J)�U3T�U��5:a��@0祚�T�6-�N�zJ��f�+�pO��(���Xv��i8�_,�"�8Yk�cY�?S����G�ș�#ޗ�M�J�s�&�������%V7�����r0��������jwQ�r�e�p�ׇ) ��Y��$�+JZ������N�V�Bv��zx��(��D��H<���yȶb?Q�S�Ԫ)� �y{n.d,d~:��K�������ŶjIMV|�0ճ��r?��G��[���i�v6"�;7	�f����Tby��Ά��tU��z6�EU�X�G?T�J�A�#�"�����25�R��-�Fy�� .Y�@���[�S�D�a|���V��y���d/�+֊_��`/!-!W�p�3�F�"͇Wo��U�(�7��G��OR� ��g��d�?T�JByT��!�'^ߑ	����lo�Z �"P�;ѯx�\`T����,��p��b��􊌷�"5'� �%6�PM1��Q\�)���;�4��J���zU�ם��e !�+RPW�d�|�0��Z!1��h��X���	� awP��{G�'�K��6����?�#�|��Û���w��h�Z���>
��7��W�f��{�k��.�I����z������pR[�����t��#�p�a�}s
l�����jæ�%2:��8?�C�ن^{/<Pn�T��z}����9Ũ`�<O���(�����b�<X`�i��2��Ko,��� �1t2��7�
@�u!�	�h�x�6�NrM�?y���4D����+;H+�(1x`z�!��	X�9���"�cmqx8F��>�Z���<F/��ؽ�E���T��pJ>!�uPD����w�q7˭B9�s�<Nb>�G/ɷ;w���� ��i����������i16\h�{F���e�'!x5��k�yG�^�T;�KC'7�P\iՋ16���o&�4,����ˏ�^r�` ��E.�{��
	�F��~^�j��J�I����*q��.���n�p��2p����7�CF/T�0�}�!���uXъ������+3��
~K�[�F!�N�$IT�˷��ĩ�-���/Ϭ�b���f�z����S_n�2J���P_\��NB���@��:�_6����[B]�=�3�s��y-����Vs�.�o-'}������c���$�[�o�,~ـ	�q�<�g�G�� rҌ$㿟.~��זV��<���,!X��|7����y�Y�	E�R��ٱ(F�mgL]2�M��哈�2z)|���@�_Z�B�ʁ�\�L������Ɯ(�׵J�=�øa�z��y赍�������a.K��{Dj���&�u���X�dl�����DDH�<�i�@���۠U��yѲ�CY^Lqg�J��/s�-�[v�R�Ā��<@8J;^�����+=ߛvľ�\xʰB�(�#V4�v��G[|15��=qˣ���tx�a3�h��80f�p��k�
�톔ګ�v��`b���2-��d��^�:N�~��/M#��ۮ�<�����>_9����D�ز�����T�#��I�� 2�g��a]>$*
"��#U�T�}n����_4��/�>UEmW���b�rx�Zf��1eyo�b��q�$ev�s�	��C�֗�W�Pl�çMS*����8%2eD�����>�L����>�y�{��Vk���srG-v�����3P��˒�gnZ}���߄�{�Tz�~��UHmj��
��7�Σ���җ9Գ��oȂ���lY�<M��9����j��n/Lc�0y���b5T�M���o!�Q֊>>�Z18�Z~^���X�a�q�uܼjV���JP���R����E��^۰M����@(M~P�7ZoY�������O�3�1*T��n�p��i�[�4��Kz�f�I��Ͽ���?��g�\΍ ���{DfQ��P�6v�J=͢�6l˅�v�C,N1}l��u(Aw`��r�� �̎���9Oǆ�H�'�G�L�j=BQ����ύ�O ��G���Sܐna�����.�"�r���.e���nIk'���׵��fY'�5^&M:���Y	2-p�`'����.�aG�iy�!I(�7g���t�;�P)쩃v�ns.��������1hn9�<����1��l�=�(�9��9��T�j�r���/�Jo=�o��7����?�(f�ǳR[k)��k�n�M���ỷ-i�ݽ)R�a1A��������O�F�m/�_Z�8{Q9��O<�-���V�V�z���c|F�	���y6ٶM���`5?̉D�P��HF�5��( ��KE���z@���x���b?��W|_jl`�?��(��W�����_�ߑ��L[�rF$"A��A$ ���k�H�����&o�um?,y&w���'��N�W;��b�|�X��JXڜ�'�5��O��g�22s�Q��sj߁o�<z)Y�u�ʦ�"H_v��R��*=���hT�Β��2��MWC���¶q�V��8�~��$��-Mr�4�A�1&S�
��n��d��)�i���Q�H�,昙�������M�����9��<���/b�F�ӦS�����O|�^���j�]����c�	ܿ3��4��X��f�.�DC'P���!0���fX�!����	�)ı�0�ر��B�V�J�m�]�e�>	D9��i�bQBKpq�t��b�恎��9�Iė<��M#j�#C���u��u�\��X�u�m)��G���Cڝn�<�1T�S�G�R6e�aэ:ӓ@�e���N����[�c)����PZ���J�i�/�K���{� h��η/� ?a�#�����A��g�5�)+-B�uMmF�"�c��#�Ҿ�J�
����vp3���Di�Ͽp��*T�C��'3�6��Ik,@:�������kS̻�.���ۅ_�.��F�3�/�aw�XlxVHYEB    fa00    12e09U�Huk������G�k~�!E[�����
��1<@O�lEi�����f�
���)�Q��n�f@�ne���kˀթp3V�!iXY��i�`�wT�|dYs8i�m�!g:Mb=�՗(��g�XʎŤf\-
�6 X�im~�&}@���'GY��v�JY�jn��!4�ߠ:k���%^-@�y<��f�\��.<�ȑEɨTmo��G�ū�E�%�y3���\�17&���|�%�n�k&�;��鼥^��FV9��Vs�hc�U�I(�Yb�N1vťJ<]��'�mc�d��4���� %�ԇ��k
ؠ3$(��B�!��-m�ԘK�z��B���y`���Z�p���RoY�6�m�l�n���H�yػ�)|o�R�9`E�1�_y-!Y՜ˁ2Ք�w�~������C Ҙ�5?���
`6W +S�� 5lR��M-�t�u���U�M�ĭ��Ð��``��UnUϺQ�>��D:����|����^�z|9������/�4΃dU��px|ĕjV��Q��v��Dh��E���wFz䤕�W��)�$$+�7\�}��)6&��Ҧ�EYQtΘS�4�����wp`�����D�Z�u_�Ȩ��]
������o*U��x��}��Ky��wJ:��l�O1������'D�o�H׮�i��U�i0�ҡʇ<�E!�a�2g������E�!������4XOy�*q$�(���)�b4eN���&f0~���A��+x��U��I4��u5�ӓ�YW��a�f�� �V
�{����G��IT�������`��`�w׸����@��4x�0��*��v@y������89Yhg�#�Pt���I�8�Bu�>��ǹ7ݯ'8�9odX�rS�ߎb|z�: �tf�*�`�n�������K�g�]�@b-�5;Ɯ�C�l��,:��*��W��_�|�V�����t_��ԓK��RǄ�\%G'��n�.����F��mǖ�V�G1B�"�i�#E�&q�[$���2s}`��0��Q�z��ϵ�~9hs"�;��{�{��>OY��h�j�����Xp�$���T8ӱ�3�7e�O��b*�D��L��}>!� <�Ύc�Y��v-���W���
��T"j��Ί�,�
�c�5Ag�)x�~5���W��ܵ�t7oMQ=�T���/��*�at0�nR2 �Q�rCg�P���	��֕ٯ2Y���Z:u��<�����e-��!�	y-P�h�^y�$�E\���O�a����R���'Z2FNs'������Z�\��B�؄F��H��՚_���g�����[d�v��'X��$����^�� ������s�-�]���i���L^����j�J�H(�Z��|�!�����T���G����*>�jq7N�L�:;;�Мݑo^�/[#�}�ٮ4/�=b�P�(�<8�SȞ@����҅��++���pǉ����{"��\D��B�<  �b<�f�[��'�5�s����ڷ������~��FYȾ[��fr���Ny����H72\_�8���y�"��
��kf"���^����M�?:>�v�H�Pe��[)�%���Lw���$-�؈V���u�8:���Y��H�Tr_����*�9H�V�j�����S@8��*��7��_���/�\��\$��q���%e�e8/+�e��GD,j\r�/*�i}�؅�_e�-�07;�M�����vl��7d�h�W�U��7k�D0�G�����������7���7�ۋ�م�N��W*5(����O��H�ז�ȭ�[�bZL�1�l�bV���W�����C�n'��%�6ܮ���3�/
����`ŷ�=$G�Q� d�Į�(��y(D$Ӄ %��,h��խQ�M�
,I��� ��i&��./~8>��s�&�*��+�vvl�X���'m��!;�����U���U �4,��>�F�_�Ņ{I@X"��!x�Kf�r�ˉ��֑��B]�*�f5�|Ȼ/K��x���k�^��C*��d�����e�X���λ����H��� ��%��ي�uGE.a2��q�����F �8i�d 7@���W�Տ���Df�˧�d��
}kTl�����;I)F�2^����1�؏j�<�@$��VzR��aa�ɤu`L����4�-�1c�����)rW�Ԟ� <����~�O������Xj�ŧ�M���$\~��O�^�={�9^7衕��-#�ҏ��{#�kՓ>��bn���#��يֳ#��p$� W�~*zR,v�(���b�S��o�j��.��$��M$�?[&����r"����U�����Q��F^��D���#�̑���u |w-h�x�)/А�O�t�"o\@��(���J���e6Tȸ�4|U�Rb$~�.ݔ�)��g����m|Y}Y'|�(�������o�t�|ܒާ��2���+�g�c�j�FH����N��K�WZ����|��c�!1��K�5��S�m��n�f�
٬��S�bW�˯�j���^�>���^(����4�1�ìe����r�7C'eEK��G|�L��G�,�ʞ�!�v�R��=w3�2}#�O2�CJ_��m���FDwn��i3.^|�{����x#]��W޺B�/L������a"�[[�",�ѻ���g�(����=\��۟�����.E�5��C�BepS��Hw��F9�ؽ�Y� I'(���S�n�����C���6�,�*�幦��턖�ѿMX���L����k�nN��lǙ-�ȍ@]�VG�K ��X�dz�Q�����EC�Q��4�Iw�Й,�_ʻ��٦��0��dǎkz�d�
���W͘ld�#�5�tY6ޮ�~:zҹx̐<�7����O�ay��b���`�y�`=�o�I>������D�F�cv׃_���>�YTW��z>F�����^.��$�|?��o��Xrf�Y�5�]�R�>V��6[�	����a�'u�GͲ�WU�,��r������tt��V�^��ua<蕢�N��"w�I�=*P\��et�ɠp}�o��`�3zd�1�§�F�(��byCX\�@�dP� s����+˙_B'
��P�v�a�t ��Z`GL�v��o-흸������:_�'�.�r?{�ǀ�J ���$� ���4p�:��>{>mc~�ᮼ�s�i<�>��!�op4���pF��L���F^�HS�=�0u۞~`���2�*>U��/&Ա,Qs�cM �i&xoWy�r��t�݌�
�J|)��?���_��tjı�qߖ|�#T^Wwk�I����`]_~9��1ʞ~�w~޲��`�^"P�A3=��8+BҲ�����U�����H/&�=�Z��8k��\0Y>��h��1�=�����$u9J�I.[�W..xq�a�z�Q�最@�~������
��!��E:�*\(�����~n��\�	�G�$%Βi��oi)�Ě4��;�c���A+�[6��tV�,V�I���rӴ8��t��9\�<�s�k㾐x�l@Q���z C2�P����T�JΪݪ��~4B�?���yv���	H���Ix����ӑ�K��>�$=ְY�vu�����n~�==ˋR�\��s4�) �ypc�l6�Ī�pm
0�9��P4�j"Y����Q]]k�l�ְ�%��_��n��+� ���D�*�����I��蹀H�l _̘5�F_xΒ�K�Xj#�l�X�����=aZ�xe�J(r�⇪���80����K��E�֓@��f
�(-(G�H�7�w�4R+�-pv���0�=�K�S�p�M���b����u^�)9��Q��YԦձ�kj������������#�ūdt$�����ӗxjX�G P�MY4&�O��<Hs��E.Co�ʄ;e���,��/p	}�=Y>���3�A��B��J}ҍ���o�//`T�Q������adx���;n�v���P�'�jk�� .ˋ��?�氏>�G��+�I���U
Ly�Jj$�g��/32�T?9�.H�pN��'��#e#9�Y�m�R����a�&�wFA�NL~ac{[v�g'J0�����HM@`r��;�й ��#��U��/������ʉ���+[aB&	���2���7��)��y���N���:�$Z��k�/GDA.Ý��"���Á�d��_�-h�fŃy�,h�F_� ��!e�{��[C�,-� 숁x��
O���>rB�� ��@7YJ�)�5�퍰����b��١��H���*�O���_פp��Q� �Pd�J~����C�*��q�Ҝhܮ`����t���ƫ�P��W�D�ٴ����+��D�;�7��b�d1�~Tۉ��N_���E�t�@��o�e&9_�c%���x.��P�BG+�:V188D�:��2�):i}��t��?!���ad��ή'��7e��{1��5�1yȢ~Lp.�C�KI�?i�����ʇFHiQ�(���*mb�-�ǡ,�:J�K�Nsؔ�$q���߃~vAPHi�@c5� e�:��j��J�����%�k	Y�F��Q�ٸ�-�ё�ݑ������O��HlL���}XZap?G�j3�>�Ĝz������s�N#�F��̀�3 z+��x9�`K;��)::���e]��F+ʩb��n�@6f�H�w��!O�}M��T�P���"]x鼍��ȑ�]���K���K�X��XlxVHYEB    fa00     f50㉧�~�U�L��E�����=t�e�A#��P#E�%�|����΀9T���ϔ�$��?-�ߥwݺϭXw�1����Z%Oڟ�])U�0&Myb?@'w�bp{oX���F��B:�hg(W�6u���l���]�3ΣU`'� Y��X�[j�w4�+�n��1
?�o��yW| ����P6'�-٘�6ُ*e�d~�)6ķ��I*�~�q��f�A����+����[��A��	�l���}��Ӱ�@o���~I���"]G޾���{�S2!�-��i�1�FaN��1�Si8���b��@������*�>�9��9b�1�tS�Z�	�C!1��ӝ��:�Th�l��)�k#!�e.�,�<���d��]���Y��Yx���#y2������^���i��;r*۱��C�rP�$��帎�f>̨�<az�����GW�g#��>V�l�� 8g�p��N�m^T�l;--���P���FD�0A�a�M�pH:=Z������/PƬ�W��S�������r�-��4R��E���E�)��y�2��< \Q��5�= ��@k�g#1ի  8��x2tsá#<e�eΨ�B��b!��V F�_��xxS1����@+��?rG��fFf�f��e�J��g�ZbKS��r�"F>�'-}��dd�����J�0sV[�AG\r[--�tۤ�Q�5�Յd��b	���aQ���D��d귡��/�x��(<"J�S��4�7Yd�����k(�`�khW��Y�C�|;�(P��h�)���"�m�/ �Jވ�d^�F��.'�t�wݡ)  "@#���
�Z)���j?�l�i!��
�n��'`֜�.����ٛ}qf���+۔��m#;P��40h����'������!��p|�'�v��L�FM�%�&t����.�h����\;ƪܡQ�1*1�ZrWF\�iA��6�.]`��$}#&"ߐ�
L?V/�G��k�B$D7� ��{��[�ǸT��[:��9��R����������E�@W\�fd2h���{�a�Lv��0��̂�pü�`��cY=�!)���GP��0���K�� ܈�zr��2�?�U	%'uy���L�$æ�/��1U��DK|����N���4V��&���� ��z�G��1��E�z�t�K��l����^!���Ї5MI�.�pq�A�KUd����FU�{�P�mc��"��c-�{ *�	���B�ւ0ApEC0x}UJc�=���_ � �pi�BcB�	��wU<
`�cyg'5}؏�N�=�����Z�Z���.�]��o�L��oee��#G����ཤ�m�(���
d�\w_z���F1r��C*�tn�4ɏ�gw�	�p���PS)�]�)<��9p���[PU�%<��%�n�4�PA�5!Q�,�i�˦j���	d��)v5-��K��t�b7OU:ފ^O�}Xt���hQ!��)6�pe�w[�8%<��0+��:�1=CS��,�R{���U*H�NDV�ı�����������gKz��pU�~c�H��2��yA���k<�V�΀B�3�8�2�`]z|�dymFH��
�����Q���1��S�G>h'O����b�9K;�uq�$5ep�V/��;\(�� J�`���筄��h��� iR�ì30J��:�������?F�i�C�=�Β́��͒ N��gGn4nH%�˛C�@�;�P��;�	M�h/25_}�����g������u�k�N���l>�����D�3x!?Dߟq�M�-�Na�'�Děb���CՌ����!iԉ&��ϊiӥ	��Z��:�C���.<�P0+y�dc*2�E�7����N�H3p�m�$f�e�PHJ�[��,.�<ċh �uH�cg#���1ub�LG�7��&����Nqj*���ѩ��S��qJVծ��{���v--�O	ݦ6�%�J�-��s�8TZ�׽�u�Y�yJ�����&�z;U����k�3e�RF^��-5L3�L���I���fh���gg�����H��� Ճ�q������̮n��Nä"��,콲ɖО�y_��ܜg����~m���l)($"R*4��v�Ar6j��J�lh���Wt[w��1�Slz��j��<�Y�f�?/A6]�$���z�7��EA�@P�!#���~2�D4?Nt1������m��)Y @(�����8$����$�a�񄉡��7p�%����P� �@7Yc����\���ZS�[�SPl�E�O����MϞ>Q#�)��W��+R�Mj����E�'Y��K�Y��Ś~�CԬ�H�3y�����!g"彏���r,8!�����D���W6B.�
��t�'Z
�)4�P�<x���[T��]�ʹ:F:v>��;�����lޣ"��Lª����(LyGd�v�k&���[�Z�:o@jԮ
�ќ�������C9Aqk:�@���S5.	�h����HFY�-+�o0|��ā�h2�5�Fr����_���Bil=Aj����%``FPp���M�ihk�w�h�B�B{�F�� ��paXo�G���QPqYD�i%]l��/b��]Y����r� w2A��/��I(:՛+/`�`ph �^�6x�C��7t!�v���4�-����'4N���eut�ǙƲ�����1ȤxI\޲w�^�L%R���h�S�Le>�)�v#����|��a�\x>J�UX1��z:�S�49�m��?��`Ɇ_��P�� ��:��x p�ωh1���2\?�������%U�EPf2j�.%�m��B�D<����?&�&	E��d��C;nu�[Ǵng�8Z�n\�(���״bR'Ŕb���\��z\�ħ3�qeC���;����.��C���t�-
�Ob��@`���h�7gԿ����^T	��K�.�%��2�a
��T������4`�e��;ן#xqۣ�҂��9+�5�M�<�&���>1P� �����덄������Ko�|�v��Ul���C4^%DP�0
s�:����J�j�
QWR��MYN�r	ȿ�����m�8xd:��C�hGH�>��8���D#�unA��1�[~�O�h�%��̞(0Y䄞O�1�#��b]MX��ʄ�O� Χ�
���C����DS�3�R��h��Mdv[��[p��d7!��?��0��ʛ&C�Z+�������~7��K�z�;|����Jr�y`����61��Rn-	#L�JϿ�ᐳC<g}Xm�1�C�3���<���N楔��3��Pbp�l��@6ǳ�c �{@?�X#j30	L~�b����M��M�b' ֛������F�"=v�����T�n]P+�����E����IԹ�ptF��p�|7�د�UOHX���_8zF�g���BZ1���o,">�u]��>Ne^��WN?�$�.G�G�|/f �����O=`�4�m��P��hT�@��cj��k�j2�h�[Z����N����Q�3_.I���/����HֆF��<��j6�'b�A�9���2C�^�cC)O�bƠj�B���IC>�¼}�����{��c��s�=݇P��uSQ��*cg�_���L�-��W����8�g�$X�N���zD����6BM?PuKN<[���J�q�"�����~u�1@0�z��<�Jv�I6���9����_�I���2ȣү)`Oa�C��8���ЯA�:�<	V�@|�]leI'�]�h]ʽZ'��ȩ�{W�Ŗ�5�}=�����3
|"]��r���p$ye��R �#ZVd�A��*�Ұ��@gC.�o�:a��d��ҧ[�P�+m��.�o��.�TgT�5S�1-gi���6�1��zJ�L1q���h����3XsKC�d�XlxVHYEB    7273     560�w�6�b�іj<��/�����O\��Ū��8�W�����ry�P�@�y��O�& ���U7��w2POGu�ݩ�[�%����g����PZq�p4�,aXz�}|j�LsH?��VV�k�}Y�ӛ���A(5w�@��s �#^:������o����ќgy
[�+� K���9΄7|�{dO8-��O�?���+�p Pj�B��@y��u�sbN�wo
��S�t�s�/b'Y�FI�`T�P����N&���
��<���X{����U/m4�!����
����l�� �	� K�
@��q����X�&b�6ly�X�J8v����V�N8b�_nw~��C�*����/�34�V�Q����t��q������U|���,V��۰ظ�(���+���r���;ۑ�b��ҏF
R�)&��ĕ�ظÞ�K������2�&���
I_�{��td �4��[%�����
-3�����̢�u�(��T@'��zS�S�%<]�o��C�+��0�k2��Ѝ:�η�|_-�`ðLh^˅V�d@8ݴ�^Z�3]K�G���<W��7����TV�ת:���#����ƌ��O�ٗ��H�GҮe�l��.�׷�gQs��E�qE/^��ώ>%'���-)���:���I�;Y=������� ���>��Hf���_t,4O��M��}6\'Uu5ݯ����x�������oq�/-)��\���k&��(YW�t�?����v��7{�13mX�II��2(n&ǖ1а���ne�
��|��{�mc���G���G��hVcmv[!K�g�bQ�� {�bV-��'����� =04x��݅9�XV~�P��>T@f�$���i���儽{i�%[ݜp���"h{'�J���[YF�!� xn���*���_�{��k��woۃ�41yU���g
�')
����`/�<|�2mSh��>U�٣��]/<�	s��F+H�,'���b`���JS�O�؉&8�j��7Ie�vSFu�3,p��H�I���cC��G�d	����������%�����=���ڞ&K"��ahG�Ι��	��&U��Q�g�r�~)��B��aMs�Z�h_X0/^"x*�5I�;z!����`�r�o�Η�`�iz���D���өU�f�1�q0I�
��Q��?���:?C�Í�i�L��&`p�qi6LS�"M��������H�8�.��8�h?�أ�7�e0�݈������ᯏU0�Ʌͱ����}	����j�������J&'�%
�R$��?����֌OiT��{}C|t�Z�Ad��(xE�